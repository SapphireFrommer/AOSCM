

module MidGap_DGWCLK (DGWClkLeftNet, DGWClkRightNet, E, SE, clk);

	//ports
	output [255:0] DGWClkRightNet;
	input SE;
	input [255:0] E;
	input clk;
	output [255:0] DGWClkLeftNet;

	//wires
	wire [255:0] DGWClkRightNet;
	wire SE;
	wire [255:0] E;
	wire [255:0] ECK;
	wire clk;
	wire [255:0] DGWClkLeftNet;

	//instances
	PREICG_X0P5B_A12TR DGWCLK_gate_0(.CK(clk), .E(E[0]), .ECK(ECK[0]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_1(.CK(clk), .E(E[1]), .ECK(ECK[1]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_10(.CK(clk), .E(E[10]), .ECK(ECK[10]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_100(.CK(clk), .E(E[100]), .ECK(ECK[100]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_101(.CK(clk), .E(E[101]), .ECK(ECK[101]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_102(.CK(clk), .E(E[102]), .ECK(ECK[102]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_103(.CK(clk), .E(E[103]), .ECK(ECK[103]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_104(.CK(clk), .E(E[104]), .ECK(ECK[104]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_105(.CK(clk), .E(E[105]), .ECK(ECK[105]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_106(.CK(clk), .E(E[106]), .ECK(ECK[106]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_107(.CK(clk), .E(E[107]), .ECK(ECK[107]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_108(.CK(clk), .E(E[108]), .ECK(ECK[108]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_109(.CK(clk), .E(E[109]), .ECK(ECK[109]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_11(.CK(clk), .E(E[11]), .ECK(ECK[11]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_110(.CK(clk), .E(E[110]), .ECK(ECK[110]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_111(.CK(clk), .E(E[111]), .ECK(ECK[111]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_112(.CK(clk), .E(E[112]), .ECK(ECK[112]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_113(.CK(clk), .E(E[113]), .ECK(ECK[113]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_114(.CK(clk), .E(E[114]), .ECK(ECK[114]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_115(.CK(clk), .E(E[115]), .ECK(ECK[115]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_116(.CK(clk), .E(E[116]), .ECK(ECK[116]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_117(.CK(clk), .E(E[117]), .ECK(ECK[117]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_118(.CK(clk), .E(E[118]), .ECK(ECK[118]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_119(.CK(clk), .E(E[119]), .ECK(ECK[119]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_12(.CK(clk), .E(E[12]), .ECK(ECK[12]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_120(.CK(clk), .E(E[120]), .ECK(ECK[120]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_121(.CK(clk), .E(E[121]), .ECK(ECK[121]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_122(.CK(clk), .E(E[122]), .ECK(ECK[122]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_123(.CK(clk), .E(E[123]), .ECK(ECK[123]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_124(.CK(clk), .E(E[124]), .ECK(ECK[124]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_125(.CK(clk), .E(E[125]), .ECK(ECK[125]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_126(.CK(clk), .E(E[126]), .ECK(ECK[126]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_127(.CK(clk), .E(E[127]), .ECK(ECK[127]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_128(.CK(clk), .E(E[128]), .ECK(ECK[128]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_129(.CK(clk), .E(E[129]), .ECK(ECK[129]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_13(.CK(clk), .E(E[13]), .ECK(ECK[13]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_130(.CK(clk), .E(E[130]), .ECK(ECK[130]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_131(.CK(clk), .E(E[131]), .ECK(ECK[131]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_132(.CK(clk), .E(E[132]), .ECK(ECK[132]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_133(.CK(clk), .E(E[133]), .ECK(ECK[133]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_134(.CK(clk), .E(E[134]), .ECK(ECK[134]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_135(.CK(clk), .E(E[135]), .ECK(ECK[135]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_136(.CK(clk), .E(E[136]), .ECK(ECK[136]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_137(.CK(clk), .E(E[137]), .ECK(ECK[137]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_138(.CK(clk), .E(E[138]), .ECK(ECK[138]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_139(.CK(clk), .E(E[139]), .ECK(ECK[139]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_14(.CK(clk), .E(E[14]), .ECK(ECK[14]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_140(.CK(clk), .E(E[140]), .ECK(ECK[140]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_141(.CK(clk), .E(E[141]), .ECK(ECK[141]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_142(.CK(clk), .E(E[142]), .ECK(ECK[142]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_143(.CK(clk), .E(E[143]), .ECK(ECK[143]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_144(.CK(clk), .E(E[144]), .ECK(ECK[144]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_145(.CK(clk), .E(E[145]), .ECK(ECK[145]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_146(.CK(clk), .E(E[146]), .ECK(ECK[146]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_147(.CK(clk), .E(E[147]), .ECK(ECK[147]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_148(.CK(clk), .E(E[148]), .ECK(ECK[148]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_149(.CK(clk), .E(E[149]), .ECK(ECK[149]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_15(.CK(clk), .E(E[15]), .ECK(ECK[15]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_150(.CK(clk), .E(E[150]), .ECK(ECK[150]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_151(.CK(clk), .E(E[151]), .ECK(ECK[151]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_152(.CK(clk), .E(E[152]), .ECK(ECK[152]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_153(.CK(clk), .E(E[153]), .ECK(ECK[153]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_154(.CK(clk), .E(E[154]), .ECK(ECK[154]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_155(.CK(clk), .E(E[155]), .ECK(ECK[155]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_156(.CK(clk), .E(E[156]), .ECK(ECK[156]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_157(.CK(clk), .E(E[157]), .ECK(ECK[157]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_158(.CK(clk), .E(E[158]), .ECK(ECK[158]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_159(.CK(clk), .E(E[159]), .ECK(ECK[159]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_16(.CK(clk), .E(E[16]), .ECK(ECK[16]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_160(.CK(clk), .E(E[160]), .ECK(ECK[160]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_161(.CK(clk), .E(E[161]), .ECK(ECK[161]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_162(.CK(clk), .E(E[162]), .ECK(ECK[162]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_163(.CK(clk), .E(E[163]), .ECK(ECK[163]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_164(.CK(clk), .E(E[164]), .ECK(ECK[164]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_165(.CK(clk), .E(E[165]), .ECK(ECK[165]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_166(.CK(clk), .E(E[166]), .ECK(ECK[166]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_167(.CK(clk), .E(E[167]), .ECK(ECK[167]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_168(.CK(clk), .E(E[168]), .ECK(ECK[168]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_169(.CK(clk), .E(E[169]), .ECK(ECK[169]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_17(.CK(clk), .E(E[17]), .ECK(ECK[17]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_170(.CK(clk), .E(E[170]), .ECK(ECK[170]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_171(.CK(clk), .E(E[171]), .ECK(ECK[171]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_172(.CK(clk), .E(E[172]), .ECK(ECK[172]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_173(.CK(clk), .E(E[173]), .ECK(ECK[173]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_174(.CK(clk), .E(E[174]), .ECK(ECK[174]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_175(.CK(clk), .E(E[175]), .ECK(ECK[175]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_176(.CK(clk), .E(E[176]), .ECK(ECK[176]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_177(.CK(clk), .E(E[177]), .ECK(ECK[177]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_178(.CK(clk), .E(E[178]), .ECK(ECK[178]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_179(.CK(clk), .E(E[179]), .ECK(ECK[179]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_18(.CK(clk), .E(E[18]), .ECK(ECK[18]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_180(.CK(clk), .E(E[180]), .ECK(ECK[180]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_181(.CK(clk), .E(E[181]), .ECK(ECK[181]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_182(.CK(clk), .E(E[182]), .ECK(ECK[182]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_183(.CK(clk), .E(E[183]), .ECK(ECK[183]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_184(.CK(clk), .E(E[184]), .ECK(ECK[184]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_185(.CK(clk), .E(E[185]), .ECK(ECK[185]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_186(.CK(clk), .E(E[186]), .ECK(ECK[186]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_187(.CK(clk), .E(E[187]), .ECK(ECK[187]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_188(.CK(clk), .E(E[188]), .ECK(ECK[188]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_189(.CK(clk), .E(E[189]), .ECK(ECK[189]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_19(.CK(clk), .E(E[19]), .ECK(ECK[19]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_190(.CK(clk), .E(E[190]), .ECK(ECK[190]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_191(.CK(clk), .E(E[191]), .ECK(ECK[191]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_192(.CK(clk), .E(E[192]), .ECK(ECK[192]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_193(.CK(clk), .E(E[193]), .ECK(ECK[193]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_194(.CK(clk), .E(E[194]), .ECK(ECK[194]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_195(.CK(clk), .E(E[195]), .ECK(ECK[195]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_196(.CK(clk), .E(E[196]), .ECK(ECK[196]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_197(.CK(clk), .E(E[197]), .ECK(ECK[197]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_198(.CK(clk), .E(E[198]), .ECK(ECK[198]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_199(.CK(clk), .E(E[199]), .ECK(ECK[199]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_2(.CK(clk), .E(E[2]), .ECK(ECK[2]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_20(.CK(clk), .E(E[20]), .ECK(ECK[20]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_200(.CK(clk), .E(E[200]), .ECK(ECK[200]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_201(.CK(clk), .E(E[201]), .ECK(ECK[201]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_202(.CK(clk), .E(E[202]), .ECK(ECK[202]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_203(.CK(clk), .E(E[203]), .ECK(ECK[203]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_204(.CK(clk), .E(E[204]), .ECK(ECK[204]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_205(.CK(clk), .E(E[205]), .ECK(ECK[205]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_206(.CK(clk), .E(E[206]), .ECK(ECK[206]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_207(.CK(clk), .E(E[207]), .ECK(ECK[207]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_208(.CK(clk), .E(E[208]), .ECK(ECK[208]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_209(.CK(clk), .E(E[209]), .ECK(ECK[209]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_21(.CK(clk), .E(E[21]), .ECK(ECK[21]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_210(.CK(clk), .E(E[210]), .ECK(ECK[210]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_211(.CK(clk), .E(E[211]), .ECK(ECK[211]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_212(.CK(clk), .E(E[212]), .ECK(ECK[212]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_213(.CK(clk), .E(E[213]), .ECK(ECK[213]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_214(.CK(clk), .E(E[214]), .ECK(ECK[214]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_215(.CK(clk), .E(E[215]), .ECK(ECK[215]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_216(.CK(clk), .E(E[216]), .ECK(ECK[216]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_217(.CK(clk), .E(E[217]), .ECK(ECK[217]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_218(.CK(clk), .E(E[218]), .ECK(ECK[218]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_219(.CK(clk), .E(E[219]), .ECK(ECK[219]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_22(.CK(clk), .E(E[22]), .ECK(ECK[22]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_220(.CK(clk), .E(E[220]), .ECK(ECK[220]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_221(.CK(clk), .E(E[221]), .ECK(ECK[221]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_222(.CK(clk), .E(E[222]), .ECK(ECK[222]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_223(.CK(clk), .E(E[223]), .ECK(ECK[223]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_224(.CK(clk), .E(E[224]), .ECK(ECK[224]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_225(.CK(clk), .E(E[225]), .ECK(ECK[225]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_226(.CK(clk), .E(E[226]), .ECK(ECK[226]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_227(.CK(clk), .E(E[227]), .ECK(ECK[227]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_228(.CK(clk), .E(E[228]), .ECK(ECK[228]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_229(.CK(clk), .E(E[229]), .ECK(ECK[229]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_23(.CK(clk), .E(E[23]), .ECK(ECK[23]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_230(.CK(clk), .E(E[230]), .ECK(ECK[230]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_231(.CK(clk), .E(E[231]), .ECK(ECK[231]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_232(.CK(clk), .E(E[232]), .ECK(ECK[232]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_233(.CK(clk), .E(E[233]), .ECK(ECK[233]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_234(.CK(clk), .E(E[234]), .ECK(ECK[234]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_235(.CK(clk), .E(E[235]), .ECK(ECK[235]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_236(.CK(clk), .E(E[236]), .ECK(ECK[236]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_237(.CK(clk), .E(E[237]), .ECK(ECK[237]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_238(.CK(clk), .E(E[238]), .ECK(ECK[238]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_239(.CK(clk), .E(E[239]), .ECK(ECK[239]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_24(.CK(clk), .E(E[24]), .ECK(ECK[24]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_240(.CK(clk), .E(E[240]), .ECK(ECK[240]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_241(.CK(clk), .E(E[241]), .ECK(ECK[241]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_242(.CK(clk), .E(E[242]), .ECK(ECK[242]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_243(.CK(clk), .E(E[243]), .ECK(ECK[243]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_244(.CK(clk), .E(E[244]), .ECK(ECK[244]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_245(.CK(clk), .E(E[245]), .ECK(ECK[245]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_246(.CK(clk), .E(E[246]), .ECK(ECK[246]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_247(.CK(clk), .E(E[247]), .ECK(ECK[247]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_248(.CK(clk), .E(E[248]), .ECK(ECK[248]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_249(.CK(clk), .E(E[249]), .ECK(ECK[249]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_25(.CK(clk), .E(E[25]), .ECK(ECK[25]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_250(.CK(clk), .E(E[250]), .ECK(ECK[250]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_251(.CK(clk), .E(E[251]), .ECK(ECK[251]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_252(.CK(clk), .E(E[252]), .ECK(ECK[252]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_253(.CK(clk), .E(E[253]), .ECK(ECK[253]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_254(.CK(clk), .E(E[254]), .ECK(ECK[254]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_255(.CK(clk), .E(E[255]), .ECK(ECK[255]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_26(.CK(clk), .E(E[26]), .ECK(ECK[26]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_27(.CK(clk), .E(E[27]), .ECK(ECK[27]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_28(.CK(clk), .E(E[28]), .ECK(ECK[28]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_29(.CK(clk), .E(E[29]), .ECK(ECK[29]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_3(.CK(clk), .E(E[3]), .ECK(ECK[3]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_30(.CK(clk), .E(E[30]), .ECK(ECK[30]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_31(.CK(clk), .E(E[31]), .ECK(ECK[31]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_32(.CK(clk), .E(E[32]), .ECK(ECK[32]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_33(.CK(clk), .E(E[33]), .ECK(ECK[33]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_34(.CK(clk), .E(E[34]), .ECK(ECK[34]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_35(.CK(clk), .E(E[35]), .ECK(ECK[35]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_36(.CK(clk), .E(E[36]), .ECK(ECK[36]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_37(.CK(clk), .E(E[37]), .ECK(ECK[37]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_38(.CK(clk), .E(E[38]), .ECK(ECK[38]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_39(.CK(clk), .E(E[39]), .ECK(ECK[39]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_4(.CK(clk), .E(E[4]), .ECK(ECK[4]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_40(.CK(clk), .E(E[40]), .ECK(ECK[40]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_41(.CK(clk), .E(E[41]), .ECK(ECK[41]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_42(.CK(clk), .E(E[42]), .ECK(ECK[42]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_43(.CK(clk), .E(E[43]), .ECK(ECK[43]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_44(.CK(clk), .E(E[44]), .ECK(ECK[44]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_45(.CK(clk), .E(E[45]), .ECK(ECK[45]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_46(.CK(clk), .E(E[46]), .ECK(ECK[46]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_47(.CK(clk), .E(E[47]), .ECK(ECK[47]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_48(.CK(clk), .E(E[48]), .ECK(ECK[48]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_49(.CK(clk), .E(E[49]), .ECK(ECK[49]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_5(.CK(clk), .E(E[5]), .ECK(ECK[5]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_50(.CK(clk), .E(E[50]), .ECK(ECK[50]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_51(.CK(clk), .E(E[51]), .ECK(ECK[51]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_52(.CK(clk), .E(E[52]), .ECK(ECK[52]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_53(.CK(clk), .E(E[53]), .ECK(ECK[53]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_54(.CK(clk), .E(E[54]), .ECK(ECK[54]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_55(.CK(clk), .E(E[55]), .ECK(ECK[55]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_56(.CK(clk), .E(E[56]), .ECK(ECK[56]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_57(.CK(clk), .E(E[57]), .ECK(ECK[57]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_58(.CK(clk), .E(E[58]), .ECK(ECK[58]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_59(.CK(clk), .E(E[59]), .ECK(ECK[59]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_6(.CK(clk), .E(E[6]), .ECK(ECK[6]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_60(.CK(clk), .E(E[60]), .ECK(ECK[60]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_61(.CK(clk), .E(E[61]), .ECK(ECK[61]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_62(.CK(clk), .E(E[62]), .ECK(ECK[62]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_63(.CK(clk), .E(E[63]), .ECK(ECK[63]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_64(.CK(clk), .E(E[64]), .ECK(ECK[64]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_65(.CK(clk), .E(E[65]), .ECK(ECK[65]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_66(.CK(clk), .E(E[66]), .ECK(ECK[66]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_67(.CK(clk), .E(E[67]), .ECK(ECK[67]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_68(.CK(clk), .E(E[68]), .ECK(ECK[68]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_69(.CK(clk), .E(E[69]), .ECK(ECK[69]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_7(.CK(clk), .E(E[7]), .ECK(ECK[7]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_70(.CK(clk), .E(E[70]), .ECK(ECK[70]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_71(.CK(clk), .E(E[71]), .ECK(ECK[71]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_72(.CK(clk), .E(E[72]), .ECK(ECK[72]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_73(.CK(clk), .E(E[73]), .ECK(ECK[73]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_74(.CK(clk), .E(E[74]), .ECK(ECK[74]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_75(.CK(clk), .E(E[75]), .ECK(ECK[75]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_76(.CK(clk), .E(E[76]), .ECK(ECK[76]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_77(.CK(clk), .E(E[77]), .ECK(ECK[77]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_78(.CK(clk), .E(E[78]), .ECK(ECK[78]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_79(.CK(clk), .E(E[79]), .ECK(ECK[79]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_8(.CK(clk), .E(E[8]), .ECK(ECK[8]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_80(.CK(clk), .E(E[80]), .ECK(ECK[80]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_81(.CK(clk), .E(E[81]), .ECK(ECK[81]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_82(.CK(clk), .E(E[82]), .ECK(ECK[82]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_83(.CK(clk), .E(E[83]), .ECK(ECK[83]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_84(.CK(clk), .E(E[84]), .ECK(ECK[84]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_85(.CK(clk), .E(E[85]), .ECK(ECK[85]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_86(.CK(clk), .E(E[86]), .ECK(ECK[86]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_87(.CK(clk), .E(E[87]), .ECK(ECK[87]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_88(.CK(clk), .E(E[88]), .ECK(ECK[88]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_89(.CK(clk), .E(E[89]), .ECK(ECK[89]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_9(.CK(clk), .E(E[9]), .ECK(ECK[9]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_90(.CK(clk), .E(E[90]), .ECK(ECK[90]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_91(.CK(clk), .E(E[91]), .ECK(ECK[91]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_92(.CK(clk), .E(E[92]), .ECK(ECK[92]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_93(.CK(clk), .E(E[93]), .ECK(ECK[93]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_94(.CK(clk), .E(E[94]), .ECK(ECK[94]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_95(.CK(clk), .E(E[95]), .ECK(ECK[95]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_96(.CK(clk), .E(E[96]), .ECK(ECK[96]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_97(.CK(clk), .E(E[97]), .ECK(ECK[97]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_98(.CK(clk), .E(E[98]), .ECK(ECK[98]), .SE(SE));
	PREICG_X0P5B_A12TR DGWCLK_gate_99(.CK(clk), .E(E[99]), .ECK(ECK[99]), .SE(SE));
	BUFH_X3M_A12TR DGWClkLeftBuff_0(.A(ECK[0]), .Y(DGWClkLeftNet[0]));
	BUFH_X3M_A12TR DGWClkLeftBuff_1(.A(ECK[1]), .Y(DGWClkLeftNet[1]));
	BUFH_X3M_A12TR DGWClkLeftBuff_10(.A(ECK[10]), .Y(DGWClkLeftNet[10]));
	BUFH_X3M_A12TR DGWClkLeftBuff_100(.A(ECK[100]), .Y(DGWClkLeftNet[100]));
	BUFH_X3M_A12TR DGWClkLeftBuff_101(.A(ECK[101]), .Y(DGWClkLeftNet[101]));
	BUFH_X3M_A12TR DGWClkLeftBuff_102(.A(ECK[102]), .Y(DGWClkLeftNet[102]));
	BUFH_X3M_A12TR DGWClkLeftBuff_103(.A(ECK[103]), .Y(DGWClkLeftNet[103]));
	BUFH_X3M_A12TR DGWClkLeftBuff_104(.A(ECK[104]), .Y(DGWClkLeftNet[104]));
	BUFH_X3M_A12TR DGWClkLeftBuff_105(.A(ECK[105]), .Y(DGWClkLeftNet[105]));
	BUFH_X3M_A12TR DGWClkLeftBuff_106(.A(ECK[106]), .Y(DGWClkLeftNet[106]));
	BUFH_X3M_A12TR DGWClkLeftBuff_107(.A(ECK[107]), .Y(DGWClkLeftNet[107]));
	BUFH_X3M_A12TR DGWClkLeftBuff_108(.A(ECK[108]), .Y(DGWClkLeftNet[108]));
	BUFH_X3M_A12TR DGWClkLeftBuff_109(.A(ECK[109]), .Y(DGWClkLeftNet[109]));
	BUFH_X3M_A12TR DGWClkLeftBuff_11(.A(ECK[11]), .Y(DGWClkLeftNet[11]));
	BUFH_X3M_A12TR DGWClkLeftBuff_110(.A(ECK[110]), .Y(DGWClkLeftNet[110]));
	BUFH_X3M_A12TR DGWClkLeftBuff_111(.A(ECK[111]), .Y(DGWClkLeftNet[111]));
	BUFH_X3M_A12TR DGWClkLeftBuff_112(.A(ECK[112]), .Y(DGWClkLeftNet[112]));
	BUFH_X3M_A12TR DGWClkLeftBuff_113(.A(ECK[113]), .Y(DGWClkLeftNet[113]));
	BUFH_X3M_A12TR DGWClkLeftBuff_114(.A(ECK[114]), .Y(DGWClkLeftNet[114]));
	BUFH_X3M_A12TR DGWClkLeftBuff_115(.A(ECK[115]), .Y(DGWClkLeftNet[115]));
	BUFH_X3M_A12TR DGWClkLeftBuff_116(.A(ECK[116]), .Y(DGWClkLeftNet[116]));
	BUFH_X3M_A12TR DGWClkLeftBuff_117(.A(ECK[117]), .Y(DGWClkLeftNet[117]));
	BUFH_X3M_A12TR DGWClkLeftBuff_118(.A(ECK[118]), .Y(DGWClkLeftNet[118]));
	BUFH_X3M_A12TR DGWClkLeftBuff_119(.A(ECK[119]), .Y(DGWClkLeftNet[119]));
	BUFH_X3M_A12TR DGWClkLeftBuff_12(.A(ECK[12]), .Y(DGWClkLeftNet[12]));
	BUFH_X3M_A12TR DGWClkLeftBuff_120(.A(ECK[120]), .Y(DGWClkLeftNet[120]));
	BUFH_X3M_A12TR DGWClkLeftBuff_121(.A(ECK[121]), .Y(DGWClkLeftNet[121]));
	BUFH_X3M_A12TR DGWClkLeftBuff_122(.A(ECK[122]), .Y(DGWClkLeftNet[122]));
	BUFH_X3M_A12TR DGWClkLeftBuff_123(.A(ECK[123]), .Y(DGWClkLeftNet[123]));
	BUFH_X3M_A12TR DGWClkLeftBuff_124(.A(ECK[124]), .Y(DGWClkLeftNet[124]));
	BUFH_X3M_A12TR DGWClkLeftBuff_125(.A(ECK[125]), .Y(DGWClkLeftNet[125]));
	BUFH_X3M_A12TR DGWClkLeftBuff_126(.A(ECK[126]), .Y(DGWClkLeftNet[126]));
	BUFH_X3M_A12TR DGWClkLeftBuff_127(.A(ECK[127]), .Y(DGWClkLeftNet[127]));
	BUFH_X3M_A12TR DGWClkLeftBuff_128(.A(ECK[128]), .Y(DGWClkLeftNet[128]));
	BUFH_X3M_A12TR DGWClkLeftBuff_129(.A(ECK[129]), .Y(DGWClkLeftNet[129]));
	BUFH_X3M_A12TR DGWClkLeftBuff_13(.A(ECK[13]), .Y(DGWClkLeftNet[13]));
	BUFH_X3M_A12TR DGWClkLeftBuff_130(.A(ECK[130]), .Y(DGWClkLeftNet[130]));
	BUFH_X3M_A12TR DGWClkLeftBuff_131(.A(ECK[131]), .Y(DGWClkLeftNet[131]));
	BUFH_X3M_A12TR DGWClkLeftBuff_132(.A(ECK[132]), .Y(DGWClkLeftNet[132]));
	BUFH_X3M_A12TR DGWClkLeftBuff_133(.A(ECK[133]), .Y(DGWClkLeftNet[133]));
	BUFH_X3M_A12TR DGWClkLeftBuff_134(.A(ECK[134]), .Y(DGWClkLeftNet[134]));
	BUFH_X3M_A12TR DGWClkLeftBuff_135(.A(ECK[135]), .Y(DGWClkLeftNet[135]));
	BUFH_X3M_A12TR DGWClkLeftBuff_136(.A(ECK[136]), .Y(DGWClkLeftNet[136]));
	BUFH_X3M_A12TR DGWClkLeftBuff_137(.A(ECK[137]), .Y(DGWClkLeftNet[137]));
	BUFH_X3M_A12TR DGWClkLeftBuff_138(.A(ECK[138]), .Y(DGWClkLeftNet[138]));
	BUFH_X3M_A12TR DGWClkLeftBuff_139(.A(ECK[139]), .Y(DGWClkLeftNet[139]));
	BUFH_X3M_A12TR DGWClkLeftBuff_14(.A(ECK[14]), .Y(DGWClkLeftNet[14]));
	BUFH_X3M_A12TR DGWClkLeftBuff_140(.A(ECK[140]), .Y(DGWClkLeftNet[140]));
	BUFH_X3M_A12TR DGWClkLeftBuff_141(.A(ECK[141]), .Y(DGWClkLeftNet[141]));
	BUFH_X3M_A12TR DGWClkLeftBuff_142(.A(ECK[142]), .Y(DGWClkLeftNet[142]));
	BUFH_X3M_A12TR DGWClkLeftBuff_143(.A(ECK[143]), .Y(DGWClkLeftNet[143]));
	BUFH_X3M_A12TR DGWClkLeftBuff_144(.A(ECK[144]), .Y(DGWClkLeftNet[144]));
	BUFH_X3M_A12TR DGWClkLeftBuff_145(.A(ECK[145]), .Y(DGWClkLeftNet[145]));
	BUFH_X3M_A12TR DGWClkLeftBuff_146(.A(ECK[146]), .Y(DGWClkLeftNet[146]));
	BUFH_X3M_A12TR DGWClkLeftBuff_147(.A(ECK[147]), .Y(DGWClkLeftNet[147]));
	BUFH_X3M_A12TR DGWClkLeftBuff_148(.A(ECK[148]), .Y(DGWClkLeftNet[148]));
	BUFH_X3M_A12TR DGWClkLeftBuff_149(.A(ECK[149]), .Y(DGWClkLeftNet[149]));
	BUFH_X3M_A12TR DGWClkLeftBuff_15(.A(ECK[15]), .Y(DGWClkLeftNet[15]));
	BUFH_X3M_A12TR DGWClkLeftBuff_150(.A(ECK[150]), .Y(DGWClkLeftNet[150]));
	BUFH_X3M_A12TR DGWClkLeftBuff_151(.A(ECK[151]), .Y(DGWClkLeftNet[151]));
	BUFH_X3M_A12TR DGWClkLeftBuff_152(.A(ECK[152]), .Y(DGWClkLeftNet[152]));
	BUFH_X3M_A12TR DGWClkLeftBuff_153(.A(ECK[153]), .Y(DGWClkLeftNet[153]));
	BUFH_X3M_A12TR DGWClkLeftBuff_154(.A(ECK[154]), .Y(DGWClkLeftNet[154]));
	BUFH_X3M_A12TR DGWClkLeftBuff_155(.A(ECK[155]), .Y(DGWClkLeftNet[155]));
	BUFH_X3M_A12TR DGWClkLeftBuff_156(.A(ECK[156]), .Y(DGWClkLeftNet[156]));
	BUFH_X3M_A12TR DGWClkLeftBuff_157(.A(ECK[157]), .Y(DGWClkLeftNet[157]));
	BUFH_X3M_A12TR DGWClkLeftBuff_158(.A(ECK[158]), .Y(DGWClkLeftNet[158]));
	BUFH_X3M_A12TR DGWClkLeftBuff_159(.A(ECK[159]), .Y(DGWClkLeftNet[159]));
	BUFH_X3M_A12TR DGWClkLeftBuff_16(.A(ECK[16]), .Y(DGWClkLeftNet[16]));
	BUFH_X3M_A12TR DGWClkLeftBuff_160(.A(ECK[160]), .Y(DGWClkLeftNet[160]));
	BUFH_X3M_A12TR DGWClkLeftBuff_161(.A(ECK[161]), .Y(DGWClkLeftNet[161]));
	BUFH_X3M_A12TR DGWClkLeftBuff_162(.A(ECK[162]), .Y(DGWClkLeftNet[162]));
	BUFH_X3M_A12TR DGWClkLeftBuff_163(.A(ECK[163]), .Y(DGWClkLeftNet[163]));
	BUFH_X3M_A12TR DGWClkLeftBuff_164(.A(ECK[164]), .Y(DGWClkLeftNet[164]));
	BUFH_X3M_A12TR DGWClkLeftBuff_165(.A(ECK[165]), .Y(DGWClkLeftNet[165]));
	BUFH_X3M_A12TR DGWClkLeftBuff_166(.A(ECK[166]), .Y(DGWClkLeftNet[166]));
	BUFH_X3M_A12TR DGWClkLeftBuff_167(.A(ECK[167]), .Y(DGWClkLeftNet[167]));
	BUFH_X3M_A12TR DGWClkLeftBuff_168(.A(ECK[168]), .Y(DGWClkLeftNet[168]));
	BUFH_X3M_A12TR DGWClkLeftBuff_169(.A(ECK[169]), .Y(DGWClkLeftNet[169]));
	BUFH_X3M_A12TR DGWClkLeftBuff_17(.A(ECK[17]), .Y(DGWClkLeftNet[17]));
	BUFH_X3M_A12TR DGWClkLeftBuff_170(.A(ECK[170]), .Y(DGWClkLeftNet[170]));
	BUFH_X3M_A12TR DGWClkLeftBuff_171(.A(ECK[171]), .Y(DGWClkLeftNet[171]));
	BUFH_X3M_A12TR DGWClkLeftBuff_172(.A(ECK[172]), .Y(DGWClkLeftNet[172]));
	BUFH_X3M_A12TR DGWClkLeftBuff_173(.A(ECK[173]), .Y(DGWClkLeftNet[173]));
	BUFH_X3M_A12TR DGWClkLeftBuff_174(.A(ECK[174]), .Y(DGWClkLeftNet[174]));
	BUFH_X3M_A12TR DGWClkLeftBuff_175(.A(ECK[175]), .Y(DGWClkLeftNet[175]));
	BUFH_X3M_A12TR DGWClkLeftBuff_176(.A(ECK[176]), .Y(DGWClkLeftNet[176]));
	BUFH_X3M_A12TR DGWClkLeftBuff_177(.A(ECK[177]), .Y(DGWClkLeftNet[177]));
	BUFH_X3M_A12TR DGWClkLeftBuff_178(.A(ECK[178]), .Y(DGWClkLeftNet[178]));
	BUFH_X3M_A12TR DGWClkLeftBuff_179(.A(ECK[179]), .Y(DGWClkLeftNet[179]));
	BUFH_X3M_A12TR DGWClkLeftBuff_18(.A(ECK[18]), .Y(DGWClkLeftNet[18]));
	BUFH_X3M_A12TR DGWClkLeftBuff_180(.A(ECK[180]), .Y(DGWClkLeftNet[180]));
	BUFH_X3M_A12TR DGWClkLeftBuff_181(.A(ECK[181]), .Y(DGWClkLeftNet[181]));
	BUFH_X3M_A12TR DGWClkLeftBuff_182(.A(ECK[182]), .Y(DGWClkLeftNet[182]));
	BUFH_X3M_A12TR DGWClkLeftBuff_183(.A(ECK[183]), .Y(DGWClkLeftNet[183]));
	BUFH_X3M_A12TR DGWClkLeftBuff_184(.A(ECK[184]), .Y(DGWClkLeftNet[184]));
	BUFH_X3M_A12TR DGWClkLeftBuff_185(.A(ECK[185]), .Y(DGWClkLeftNet[185]));
	BUFH_X3M_A12TR DGWClkLeftBuff_186(.A(ECK[186]), .Y(DGWClkLeftNet[186]));
	BUFH_X3M_A12TR DGWClkLeftBuff_187(.A(ECK[187]), .Y(DGWClkLeftNet[187]));
	BUFH_X3M_A12TR DGWClkLeftBuff_188(.A(ECK[188]), .Y(DGWClkLeftNet[188]));
	BUFH_X3M_A12TR DGWClkLeftBuff_189(.A(ECK[189]), .Y(DGWClkLeftNet[189]));
	BUFH_X3M_A12TR DGWClkLeftBuff_19(.A(ECK[19]), .Y(DGWClkLeftNet[19]));
	BUFH_X3M_A12TR DGWClkLeftBuff_190(.A(ECK[190]), .Y(DGWClkLeftNet[190]));
	BUFH_X3M_A12TR DGWClkLeftBuff_191(.A(ECK[191]), .Y(DGWClkLeftNet[191]));
	BUFH_X3M_A12TR DGWClkLeftBuff_192(.A(ECK[192]), .Y(DGWClkLeftNet[192]));
	BUFH_X3M_A12TR DGWClkLeftBuff_193(.A(ECK[193]), .Y(DGWClkLeftNet[193]));
	BUFH_X3M_A12TR DGWClkLeftBuff_194(.A(ECK[194]), .Y(DGWClkLeftNet[194]));
	BUFH_X3M_A12TR DGWClkLeftBuff_195(.A(ECK[195]), .Y(DGWClkLeftNet[195]));
	BUFH_X3M_A12TR DGWClkLeftBuff_196(.A(ECK[196]), .Y(DGWClkLeftNet[196]));
	BUFH_X3M_A12TR DGWClkLeftBuff_197(.A(ECK[197]), .Y(DGWClkLeftNet[197]));
	BUFH_X3M_A12TR DGWClkLeftBuff_198(.A(ECK[198]), .Y(DGWClkLeftNet[198]));
	BUFH_X3M_A12TR DGWClkLeftBuff_199(.A(ECK[199]), .Y(DGWClkLeftNet[199]));
	BUFH_X3M_A12TR DGWClkLeftBuff_2(.A(ECK[2]), .Y(DGWClkLeftNet[2]));
	BUFH_X3M_A12TR DGWClkLeftBuff_20(.A(ECK[20]), .Y(DGWClkLeftNet[20]));
	BUFH_X3M_A12TR DGWClkLeftBuff_200(.A(ECK[200]), .Y(DGWClkLeftNet[200]));
	BUFH_X3M_A12TR DGWClkLeftBuff_201(.A(ECK[201]), .Y(DGWClkLeftNet[201]));
	BUFH_X3M_A12TR DGWClkLeftBuff_202(.A(ECK[202]), .Y(DGWClkLeftNet[202]));
	BUFH_X3M_A12TR DGWClkLeftBuff_203(.A(ECK[203]), .Y(DGWClkLeftNet[203]));
	BUFH_X3M_A12TR DGWClkLeftBuff_204(.A(ECK[204]), .Y(DGWClkLeftNet[204]));
	BUFH_X3M_A12TR DGWClkLeftBuff_205(.A(ECK[205]), .Y(DGWClkLeftNet[205]));
	BUFH_X3M_A12TR DGWClkLeftBuff_206(.A(ECK[206]), .Y(DGWClkLeftNet[206]));
	BUFH_X3M_A12TR DGWClkLeftBuff_207(.A(ECK[207]), .Y(DGWClkLeftNet[207]));
	BUFH_X3M_A12TR DGWClkLeftBuff_208(.A(ECK[208]), .Y(DGWClkLeftNet[208]));
	BUFH_X3M_A12TR DGWClkLeftBuff_209(.A(ECK[209]), .Y(DGWClkLeftNet[209]));
	BUFH_X3M_A12TR DGWClkLeftBuff_21(.A(ECK[21]), .Y(DGWClkLeftNet[21]));
	BUFH_X3M_A12TR DGWClkLeftBuff_210(.A(ECK[210]), .Y(DGWClkLeftNet[210]));
	BUFH_X3M_A12TR DGWClkLeftBuff_211(.A(ECK[211]), .Y(DGWClkLeftNet[211]));
	BUFH_X3M_A12TR DGWClkLeftBuff_212(.A(ECK[212]), .Y(DGWClkLeftNet[212]));
	BUFH_X3M_A12TR DGWClkLeftBuff_213(.A(ECK[213]), .Y(DGWClkLeftNet[213]));
	BUFH_X3M_A12TR DGWClkLeftBuff_214(.A(ECK[214]), .Y(DGWClkLeftNet[214]));
	BUFH_X3M_A12TR DGWClkLeftBuff_215(.A(ECK[215]), .Y(DGWClkLeftNet[215]));
	BUFH_X3M_A12TR DGWClkLeftBuff_216(.A(ECK[216]), .Y(DGWClkLeftNet[216]));
	BUFH_X3M_A12TR DGWClkLeftBuff_217(.A(ECK[217]), .Y(DGWClkLeftNet[217]));
	BUFH_X3M_A12TR DGWClkLeftBuff_218(.A(ECK[218]), .Y(DGWClkLeftNet[218]));
	BUFH_X3M_A12TR DGWClkLeftBuff_219(.A(ECK[219]), .Y(DGWClkLeftNet[219]));
	BUFH_X3M_A12TR DGWClkLeftBuff_22(.A(ECK[22]), .Y(DGWClkLeftNet[22]));
	BUFH_X3M_A12TR DGWClkLeftBuff_220(.A(ECK[220]), .Y(DGWClkLeftNet[220]));
	BUFH_X3M_A12TR DGWClkLeftBuff_221(.A(ECK[221]), .Y(DGWClkLeftNet[221]));
	BUFH_X3M_A12TR DGWClkLeftBuff_222(.A(ECK[222]), .Y(DGWClkLeftNet[222]));
	BUFH_X3M_A12TR DGWClkLeftBuff_223(.A(ECK[223]), .Y(DGWClkLeftNet[223]));
	BUFH_X3M_A12TR DGWClkLeftBuff_224(.A(ECK[224]), .Y(DGWClkLeftNet[224]));
	BUFH_X3M_A12TR DGWClkLeftBuff_225(.A(ECK[225]), .Y(DGWClkLeftNet[225]));
	BUFH_X3M_A12TR DGWClkLeftBuff_226(.A(ECK[226]), .Y(DGWClkLeftNet[226]));
	BUFH_X3M_A12TR DGWClkLeftBuff_227(.A(ECK[227]), .Y(DGWClkLeftNet[227]));
	BUFH_X3M_A12TR DGWClkLeftBuff_228(.A(ECK[228]), .Y(DGWClkLeftNet[228]));
	BUFH_X3M_A12TR DGWClkLeftBuff_229(.A(ECK[229]), .Y(DGWClkLeftNet[229]));
	BUFH_X3M_A12TR DGWClkLeftBuff_23(.A(ECK[23]), .Y(DGWClkLeftNet[23]));
	BUFH_X3M_A12TR DGWClkLeftBuff_230(.A(ECK[230]), .Y(DGWClkLeftNet[230]));
	BUFH_X3M_A12TR DGWClkLeftBuff_231(.A(ECK[231]), .Y(DGWClkLeftNet[231]));
	BUFH_X3M_A12TR DGWClkLeftBuff_232(.A(ECK[232]), .Y(DGWClkLeftNet[232]));
	BUFH_X3M_A12TR DGWClkLeftBuff_233(.A(ECK[233]), .Y(DGWClkLeftNet[233]));
	BUFH_X3M_A12TR DGWClkLeftBuff_234(.A(ECK[234]), .Y(DGWClkLeftNet[234]));
	BUFH_X3M_A12TR DGWClkLeftBuff_235(.A(ECK[235]), .Y(DGWClkLeftNet[235]));
	BUFH_X3M_A12TR DGWClkLeftBuff_236(.A(ECK[236]), .Y(DGWClkLeftNet[236]));
	BUFH_X3M_A12TR DGWClkLeftBuff_237(.A(ECK[237]), .Y(DGWClkLeftNet[237]));
	BUFH_X3M_A12TR DGWClkLeftBuff_238(.A(ECK[238]), .Y(DGWClkLeftNet[238]));
	BUFH_X3M_A12TR DGWClkLeftBuff_239(.A(ECK[239]), .Y(DGWClkLeftNet[239]));
	BUFH_X3M_A12TR DGWClkLeftBuff_24(.A(ECK[24]), .Y(DGWClkLeftNet[24]));
	BUFH_X3M_A12TR DGWClkLeftBuff_240(.A(ECK[240]), .Y(DGWClkLeftNet[240]));
	BUFH_X3M_A12TR DGWClkLeftBuff_241(.A(ECK[241]), .Y(DGWClkLeftNet[241]));
	BUFH_X3M_A12TR DGWClkLeftBuff_242(.A(ECK[242]), .Y(DGWClkLeftNet[242]));
	BUFH_X3M_A12TR DGWClkLeftBuff_243(.A(ECK[243]), .Y(DGWClkLeftNet[243]));
	BUFH_X3M_A12TR DGWClkLeftBuff_244(.A(ECK[244]), .Y(DGWClkLeftNet[244]));
	BUFH_X3M_A12TR DGWClkLeftBuff_245(.A(ECK[245]), .Y(DGWClkLeftNet[245]));
	BUFH_X3M_A12TR DGWClkLeftBuff_246(.A(ECK[246]), .Y(DGWClkLeftNet[246]));
	BUFH_X3M_A12TR DGWClkLeftBuff_247(.A(ECK[247]), .Y(DGWClkLeftNet[247]));
	BUFH_X3M_A12TR DGWClkLeftBuff_248(.A(ECK[248]), .Y(DGWClkLeftNet[248]));
	BUFH_X3M_A12TR DGWClkLeftBuff_249(.A(ECK[249]), .Y(DGWClkLeftNet[249]));
	BUFH_X3M_A12TR DGWClkLeftBuff_25(.A(ECK[25]), .Y(DGWClkLeftNet[25]));
	BUFH_X3M_A12TR DGWClkLeftBuff_250(.A(ECK[250]), .Y(DGWClkLeftNet[250]));
	BUFH_X3M_A12TR DGWClkLeftBuff_251(.A(ECK[251]), .Y(DGWClkLeftNet[251]));
	BUFH_X3M_A12TR DGWClkLeftBuff_252(.A(ECK[252]), .Y(DGWClkLeftNet[252]));
	BUFH_X3M_A12TR DGWClkLeftBuff_253(.A(ECK[253]), .Y(DGWClkLeftNet[253]));
	BUFH_X3M_A12TR DGWClkLeftBuff_254(.A(ECK[254]), .Y(DGWClkLeftNet[254]));
	BUFH_X3M_A12TR DGWClkLeftBuff_255(.A(ECK[255]), .Y(DGWClkLeftNet[255]));
	BUFH_X3M_A12TR DGWClkLeftBuff_26(.A(ECK[26]), .Y(DGWClkLeftNet[26]));
	BUFH_X3M_A12TR DGWClkLeftBuff_27(.A(ECK[27]), .Y(DGWClkLeftNet[27]));
	BUFH_X3M_A12TR DGWClkLeftBuff_28(.A(ECK[28]), .Y(DGWClkLeftNet[28]));
	BUFH_X3M_A12TR DGWClkLeftBuff_29(.A(ECK[29]), .Y(DGWClkLeftNet[29]));
	BUFH_X3M_A12TR DGWClkLeftBuff_3(.A(ECK[3]), .Y(DGWClkLeftNet[3]));
	BUFH_X3M_A12TR DGWClkLeftBuff_30(.A(ECK[30]), .Y(DGWClkLeftNet[30]));
	BUFH_X3M_A12TR DGWClkLeftBuff_31(.A(ECK[31]), .Y(DGWClkLeftNet[31]));
	BUFH_X3M_A12TR DGWClkLeftBuff_32(.A(ECK[32]), .Y(DGWClkLeftNet[32]));
	BUFH_X3M_A12TR DGWClkLeftBuff_33(.A(ECK[33]), .Y(DGWClkLeftNet[33]));
	BUFH_X3M_A12TR DGWClkLeftBuff_34(.A(ECK[34]), .Y(DGWClkLeftNet[34]));
	BUFH_X3M_A12TR DGWClkLeftBuff_35(.A(ECK[35]), .Y(DGWClkLeftNet[35]));
	BUFH_X3M_A12TR DGWClkLeftBuff_36(.A(ECK[36]), .Y(DGWClkLeftNet[36]));
	BUFH_X3M_A12TR DGWClkLeftBuff_37(.A(ECK[37]), .Y(DGWClkLeftNet[37]));
	BUFH_X3M_A12TR DGWClkLeftBuff_38(.A(ECK[38]), .Y(DGWClkLeftNet[38]));
	BUFH_X3M_A12TR DGWClkLeftBuff_39(.A(ECK[39]), .Y(DGWClkLeftNet[39]));
	BUFH_X3M_A12TR DGWClkLeftBuff_4(.A(ECK[4]), .Y(DGWClkLeftNet[4]));
	BUFH_X3M_A12TR DGWClkLeftBuff_40(.A(ECK[40]), .Y(DGWClkLeftNet[40]));
	BUFH_X3M_A12TR DGWClkLeftBuff_41(.A(ECK[41]), .Y(DGWClkLeftNet[41]));
	BUFH_X3M_A12TR DGWClkLeftBuff_42(.A(ECK[42]), .Y(DGWClkLeftNet[42]));
	BUFH_X3M_A12TR DGWClkLeftBuff_43(.A(ECK[43]), .Y(DGWClkLeftNet[43]));
	BUFH_X3M_A12TR DGWClkLeftBuff_44(.A(ECK[44]), .Y(DGWClkLeftNet[44]));
	BUFH_X3M_A12TR DGWClkLeftBuff_45(.A(ECK[45]), .Y(DGWClkLeftNet[45]));
	BUFH_X3M_A12TR DGWClkLeftBuff_46(.A(ECK[46]), .Y(DGWClkLeftNet[46]));
	BUFH_X3M_A12TR DGWClkLeftBuff_47(.A(ECK[47]), .Y(DGWClkLeftNet[47]));
	BUFH_X3M_A12TR DGWClkLeftBuff_48(.A(ECK[48]), .Y(DGWClkLeftNet[48]));
	BUFH_X3M_A12TR DGWClkLeftBuff_49(.A(ECK[49]), .Y(DGWClkLeftNet[49]));
	BUFH_X3M_A12TR DGWClkLeftBuff_5(.A(ECK[5]), .Y(DGWClkLeftNet[5]));
	BUFH_X3M_A12TR DGWClkLeftBuff_50(.A(ECK[50]), .Y(DGWClkLeftNet[50]));
	BUFH_X3M_A12TR DGWClkLeftBuff_51(.A(ECK[51]), .Y(DGWClkLeftNet[51]));
	BUFH_X3M_A12TR DGWClkLeftBuff_52(.A(ECK[52]), .Y(DGWClkLeftNet[52]));
	BUFH_X3M_A12TR DGWClkLeftBuff_53(.A(ECK[53]), .Y(DGWClkLeftNet[53]));
	BUFH_X3M_A12TR DGWClkLeftBuff_54(.A(ECK[54]), .Y(DGWClkLeftNet[54]));
	BUFH_X3M_A12TR DGWClkLeftBuff_55(.A(ECK[55]), .Y(DGWClkLeftNet[55]));
	BUFH_X3M_A12TR DGWClkLeftBuff_56(.A(ECK[56]), .Y(DGWClkLeftNet[56]));
	BUFH_X3M_A12TR DGWClkLeftBuff_57(.A(ECK[57]), .Y(DGWClkLeftNet[57]));
	BUFH_X3M_A12TR DGWClkLeftBuff_58(.A(ECK[58]), .Y(DGWClkLeftNet[58]));
	BUFH_X3M_A12TR DGWClkLeftBuff_59(.A(ECK[59]), .Y(DGWClkLeftNet[59]));
	BUFH_X3M_A12TR DGWClkLeftBuff_6(.A(ECK[6]), .Y(DGWClkLeftNet[6]));
	BUFH_X3M_A12TR DGWClkLeftBuff_60(.A(ECK[60]), .Y(DGWClkLeftNet[60]));
	BUFH_X3M_A12TR DGWClkLeftBuff_61(.A(ECK[61]), .Y(DGWClkLeftNet[61]));
	BUFH_X3M_A12TR DGWClkLeftBuff_62(.A(ECK[62]), .Y(DGWClkLeftNet[62]));
	BUFH_X3M_A12TR DGWClkLeftBuff_63(.A(ECK[63]), .Y(DGWClkLeftNet[63]));
	BUFH_X3M_A12TR DGWClkLeftBuff_64(.A(ECK[64]), .Y(DGWClkLeftNet[64]));
	BUFH_X3M_A12TR DGWClkLeftBuff_65(.A(ECK[65]), .Y(DGWClkLeftNet[65]));
	BUFH_X3M_A12TR DGWClkLeftBuff_66(.A(ECK[66]), .Y(DGWClkLeftNet[66]));
	BUFH_X3M_A12TR DGWClkLeftBuff_67(.A(ECK[67]), .Y(DGWClkLeftNet[67]));
	BUFH_X3M_A12TR DGWClkLeftBuff_68(.A(ECK[68]), .Y(DGWClkLeftNet[68]));
	BUFH_X3M_A12TR DGWClkLeftBuff_69(.A(ECK[69]), .Y(DGWClkLeftNet[69]));
	BUFH_X3M_A12TR DGWClkLeftBuff_7(.A(ECK[7]), .Y(DGWClkLeftNet[7]));
	BUFH_X3M_A12TR DGWClkLeftBuff_70(.A(ECK[70]), .Y(DGWClkLeftNet[70]));
	BUFH_X3M_A12TR DGWClkLeftBuff_71(.A(ECK[71]), .Y(DGWClkLeftNet[71]));
	BUFH_X3M_A12TR DGWClkLeftBuff_72(.A(ECK[72]), .Y(DGWClkLeftNet[72]));
	BUFH_X3M_A12TR DGWClkLeftBuff_73(.A(ECK[73]), .Y(DGWClkLeftNet[73]));
	BUFH_X3M_A12TR DGWClkLeftBuff_74(.A(ECK[74]), .Y(DGWClkLeftNet[74]));
	BUFH_X3M_A12TR DGWClkLeftBuff_75(.A(ECK[75]), .Y(DGWClkLeftNet[75]));
	BUFH_X3M_A12TR DGWClkLeftBuff_76(.A(ECK[76]), .Y(DGWClkLeftNet[76]));
	BUFH_X3M_A12TR DGWClkLeftBuff_77(.A(ECK[77]), .Y(DGWClkLeftNet[77]));
	BUFH_X3M_A12TR DGWClkLeftBuff_78(.A(ECK[78]), .Y(DGWClkLeftNet[78]));
	BUFH_X3M_A12TR DGWClkLeftBuff_79(.A(ECK[79]), .Y(DGWClkLeftNet[79]));
	BUFH_X3M_A12TR DGWClkLeftBuff_8(.A(ECK[8]), .Y(DGWClkLeftNet[8]));
	BUFH_X3M_A12TR DGWClkLeftBuff_80(.A(ECK[80]), .Y(DGWClkLeftNet[80]));
	BUFH_X3M_A12TR DGWClkLeftBuff_81(.A(ECK[81]), .Y(DGWClkLeftNet[81]));
	BUFH_X3M_A12TR DGWClkLeftBuff_82(.A(ECK[82]), .Y(DGWClkLeftNet[82]));
	BUFH_X3M_A12TR DGWClkLeftBuff_83(.A(ECK[83]), .Y(DGWClkLeftNet[83]));
	BUFH_X3M_A12TR DGWClkLeftBuff_84(.A(ECK[84]), .Y(DGWClkLeftNet[84]));
	BUFH_X3M_A12TR DGWClkLeftBuff_85(.A(ECK[85]), .Y(DGWClkLeftNet[85]));
	BUFH_X3M_A12TR DGWClkLeftBuff_86(.A(ECK[86]), .Y(DGWClkLeftNet[86]));
	BUFH_X3M_A12TR DGWClkLeftBuff_87(.A(ECK[87]), .Y(DGWClkLeftNet[87]));
	BUFH_X3M_A12TR DGWClkLeftBuff_88(.A(ECK[88]), .Y(DGWClkLeftNet[88]));
	BUFH_X3M_A12TR DGWClkLeftBuff_89(.A(ECK[89]), .Y(DGWClkLeftNet[89]));
	BUFH_X3M_A12TR DGWClkLeftBuff_9(.A(ECK[9]), .Y(DGWClkLeftNet[9]));
	BUFH_X3M_A12TR DGWClkLeftBuff_90(.A(ECK[90]), .Y(DGWClkLeftNet[90]));
	BUFH_X3M_A12TR DGWClkLeftBuff_91(.A(ECK[91]), .Y(DGWClkLeftNet[91]));
	BUFH_X3M_A12TR DGWClkLeftBuff_92(.A(ECK[92]), .Y(DGWClkLeftNet[92]));
	BUFH_X3M_A12TR DGWClkLeftBuff_93(.A(ECK[93]), .Y(DGWClkLeftNet[93]));
	BUFH_X3M_A12TR DGWClkLeftBuff_94(.A(ECK[94]), .Y(DGWClkLeftNet[94]));
	BUFH_X3M_A12TR DGWClkLeftBuff_95(.A(ECK[95]), .Y(DGWClkLeftNet[95]));
	BUFH_X3M_A12TR DGWClkLeftBuff_96(.A(ECK[96]), .Y(DGWClkLeftNet[96]));
	BUFH_X3M_A12TR DGWClkLeftBuff_97(.A(ECK[97]), .Y(DGWClkLeftNet[97]));
	BUFH_X3M_A12TR DGWClkLeftBuff_98(.A(ECK[98]), .Y(DGWClkLeftNet[98]));
	BUFH_X3M_A12TR DGWClkLeftBuff_99(.A(ECK[99]), .Y(DGWClkLeftNet[99]));
	BUFH_X3M_A12TR DGWClkRightBuff_0(.A(ECK[0]), .Y(DGWClkRightNet[0]));
	BUFH_X3M_A12TR DGWClkRightBuff_1(.A(ECK[1]), .Y(DGWClkRightNet[1]));
	BUFH_X3M_A12TR DGWClkRightBuff_10(.A(ECK[10]), .Y(DGWClkRightNet[10]));
	BUFH_X3M_A12TR DGWClkRightBuff_100(.A(ECK[100]), .Y(DGWClkRightNet[100]));
	BUFH_X3M_A12TR DGWClkRightBuff_101(.A(ECK[101]), .Y(DGWClkRightNet[101]));
	BUFH_X3M_A12TR DGWClkRightBuff_102(.A(ECK[102]), .Y(DGWClkRightNet[102]));
	BUFH_X3M_A12TR DGWClkRightBuff_103(.A(ECK[103]), .Y(DGWClkRightNet[103]));
	BUFH_X3M_A12TR DGWClkRightBuff_104(.A(ECK[104]), .Y(DGWClkRightNet[104]));
	BUFH_X3M_A12TR DGWClkRightBuff_105(.A(ECK[105]), .Y(DGWClkRightNet[105]));
	BUFH_X3M_A12TR DGWClkRightBuff_106(.A(ECK[106]), .Y(DGWClkRightNet[106]));
	BUFH_X3M_A12TR DGWClkRightBuff_107(.A(ECK[107]), .Y(DGWClkRightNet[107]));
	BUFH_X3M_A12TR DGWClkRightBuff_108(.A(ECK[108]), .Y(DGWClkRightNet[108]));
	BUFH_X3M_A12TR DGWClkRightBuff_109(.A(ECK[109]), .Y(DGWClkRightNet[109]));
	BUFH_X3M_A12TR DGWClkRightBuff_11(.A(ECK[11]), .Y(DGWClkRightNet[11]));
	BUFH_X3M_A12TR DGWClkRightBuff_110(.A(ECK[110]), .Y(DGWClkRightNet[110]));
	BUFH_X3M_A12TR DGWClkRightBuff_111(.A(ECK[111]), .Y(DGWClkRightNet[111]));
	BUFH_X3M_A12TR DGWClkRightBuff_112(.A(ECK[112]), .Y(DGWClkRightNet[112]));
	BUFH_X3M_A12TR DGWClkRightBuff_113(.A(ECK[113]), .Y(DGWClkRightNet[113]));
	BUFH_X3M_A12TR DGWClkRightBuff_114(.A(ECK[114]), .Y(DGWClkRightNet[114]));
	BUFH_X3M_A12TR DGWClkRightBuff_115(.A(ECK[115]), .Y(DGWClkRightNet[115]));
	BUFH_X3M_A12TR DGWClkRightBuff_116(.A(ECK[116]), .Y(DGWClkRightNet[116]));
	BUFH_X3M_A12TR DGWClkRightBuff_117(.A(ECK[117]), .Y(DGWClkRightNet[117]));
	BUFH_X3M_A12TR DGWClkRightBuff_118(.A(ECK[118]), .Y(DGWClkRightNet[118]));
	BUFH_X3M_A12TR DGWClkRightBuff_119(.A(ECK[119]), .Y(DGWClkRightNet[119]));
	BUFH_X3M_A12TR DGWClkRightBuff_12(.A(ECK[12]), .Y(DGWClkRightNet[12]));
	BUFH_X3M_A12TR DGWClkRightBuff_120(.A(ECK[120]), .Y(DGWClkRightNet[120]));
	BUFH_X3M_A12TR DGWClkRightBuff_121(.A(ECK[121]), .Y(DGWClkRightNet[121]));
	BUFH_X3M_A12TR DGWClkRightBuff_122(.A(ECK[122]), .Y(DGWClkRightNet[122]));
	BUFH_X3M_A12TR DGWClkRightBuff_123(.A(ECK[123]), .Y(DGWClkRightNet[123]));
	BUFH_X3M_A12TR DGWClkRightBuff_124(.A(ECK[124]), .Y(DGWClkRightNet[124]));
	BUFH_X3M_A12TR DGWClkRightBuff_125(.A(ECK[125]), .Y(DGWClkRightNet[125]));
	BUFH_X3M_A12TR DGWClkRightBuff_126(.A(ECK[126]), .Y(DGWClkRightNet[126]));
	BUFH_X3M_A12TR DGWClkRightBuff_127(.A(ECK[127]), .Y(DGWClkRightNet[127]));
	BUFH_X3M_A12TR DGWClkRightBuff_128(.A(ECK[128]), .Y(DGWClkRightNet[128]));
	BUFH_X3M_A12TR DGWClkRightBuff_129(.A(ECK[129]), .Y(DGWClkRightNet[129]));
	BUFH_X3M_A12TR DGWClkRightBuff_13(.A(ECK[13]), .Y(DGWClkRightNet[13]));
	BUFH_X3M_A12TR DGWClkRightBuff_130(.A(ECK[130]), .Y(DGWClkRightNet[130]));
	BUFH_X3M_A12TR DGWClkRightBuff_131(.A(ECK[131]), .Y(DGWClkRightNet[131]));
	BUFH_X3M_A12TR DGWClkRightBuff_132(.A(ECK[132]), .Y(DGWClkRightNet[132]));
	BUFH_X3M_A12TR DGWClkRightBuff_133(.A(ECK[133]), .Y(DGWClkRightNet[133]));
	BUFH_X3M_A12TR DGWClkRightBuff_134(.A(ECK[134]), .Y(DGWClkRightNet[134]));
	BUFH_X3M_A12TR DGWClkRightBuff_135(.A(ECK[135]), .Y(DGWClkRightNet[135]));
	BUFH_X3M_A12TR DGWClkRightBuff_136(.A(ECK[136]), .Y(DGWClkRightNet[136]));
	BUFH_X3M_A12TR DGWClkRightBuff_137(.A(ECK[137]), .Y(DGWClkRightNet[137]));
	BUFH_X3M_A12TR DGWClkRightBuff_138(.A(ECK[138]), .Y(DGWClkRightNet[138]));
	BUFH_X3M_A12TR DGWClkRightBuff_139(.A(ECK[139]), .Y(DGWClkRightNet[139]));
	BUFH_X3M_A12TR DGWClkRightBuff_14(.A(ECK[14]), .Y(DGWClkRightNet[14]));
	BUFH_X3M_A12TR DGWClkRightBuff_140(.A(ECK[140]), .Y(DGWClkRightNet[140]));
	BUFH_X3M_A12TR DGWClkRightBuff_141(.A(ECK[141]), .Y(DGWClkRightNet[141]));
	BUFH_X3M_A12TR DGWClkRightBuff_142(.A(ECK[142]), .Y(DGWClkRightNet[142]));
	BUFH_X3M_A12TR DGWClkRightBuff_143(.A(ECK[143]), .Y(DGWClkRightNet[143]));
	BUFH_X3M_A12TR DGWClkRightBuff_144(.A(ECK[144]), .Y(DGWClkRightNet[144]));
	BUFH_X3M_A12TR DGWClkRightBuff_145(.A(ECK[145]), .Y(DGWClkRightNet[145]));
	BUFH_X3M_A12TR DGWClkRightBuff_146(.A(ECK[146]), .Y(DGWClkRightNet[146]));
	BUFH_X3M_A12TR DGWClkRightBuff_147(.A(ECK[147]), .Y(DGWClkRightNet[147]));
	BUFH_X3M_A12TR DGWClkRightBuff_148(.A(ECK[148]), .Y(DGWClkRightNet[148]));
	BUFH_X3M_A12TR DGWClkRightBuff_149(.A(ECK[149]), .Y(DGWClkRightNet[149]));
	BUFH_X3M_A12TR DGWClkRightBuff_15(.A(ECK[15]), .Y(DGWClkRightNet[15]));
	BUFH_X3M_A12TR DGWClkRightBuff_150(.A(ECK[150]), .Y(DGWClkRightNet[150]));
	BUFH_X3M_A12TR DGWClkRightBuff_151(.A(ECK[151]), .Y(DGWClkRightNet[151]));
	BUFH_X3M_A12TR DGWClkRightBuff_152(.A(ECK[152]), .Y(DGWClkRightNet[152]));
	BUFH_X3M_A12TR DGWClkRightBuff_153(.A(ECK[153]), .Y(DGWClkRightNet[153]));
	BUFH_X3M_A12TR DGWClkRightBuff_154(.A(ECK[154]), .Y(DGWClkRightNet[154]));
	BUFH_X3M_A12TR DGWClkRightBuff_155(.A(ECK[155]), .Y(DGWClkRightNet[155]));
	BUFH_X3M_A12TR DGWClkRightBuff_156(.A(ECK[156]), .Y(DGWClkRightNet[156]));
	BUFH_X3M_A12TR DGWClkRightBuff_157(.A(ECK[157]), .Y(DGWClkRightNet[157]));
	BUFH_X3M_A12TR DGWClkRightBuff_158(.A(ECK[158]), .Y(DGWClkRightNet[158]));
	BUFH_X3M_A12TR DGWClkRightBuff_159(.A(ECK[159]), .Y(DGWClkRightNet[159]));
	BUFH_X3M_A12TR DGWClkRightBuff_16(.A(ECK[16]), .Y(DGWClkRightNet[16]));
	BUFH_X3M_A12TR DGWClkRightBuff_160(.A(ECK[160]), .Y(DGWClkRightNet[160]));
	BUFH_X3M_A12TR DGWClkRightBuff_161(.A(ECK[161]), .Y(DGWClkRightNet[161]));
	BUFH_X3M_A12TR DGWClkRightBuff_162(.A(ECK[162]), .Y(DGWClkRightNet[162]));
	BUFH_X3M_A12TR DGWClkRightBuff_163(.A(ECK[163]), .Y(DGWClkRightNet[163]));
	BUFH_X3M_A12TR DGWClkRightBuff_164(.A(ECK[164]), .Y(DGWClkRightNet[164]));
	BUFH_X3M_A12TR DGWClkRightBuff_165(.A(ECK[165]), .Y(DGWClkRightNet[165]));
	BUFH_X3M_A12TR DGWClkRightBuff_166(.A(ECK[166]), .Y(DGWClkRightNet[166]));
	BUFH_X3M_A12TR DGWClkRightBuff_167(.A(ECK[167]), .Y(DGWClkRightNet[167]));
	BUFH_X3M_A12TR DGWClkRightBuff_168(.A(ECK[168]), .Y(DGWClkRightNet[168]));
	BUFH_X3M_A12TR DGWClkRightBuff_169(.A(ECK[169]), .Y(DGWClkRightNet[169]));
	BUFH_X3M_A12TR DGWClkRightBuff_17(.A(ECK[17]), .Y(DGWClkRightNet[17]));
	BUFH_X3M_A12TR DGWClkRightBuff_170(.A(ECK[170]), .Y(DGWClkRightNet[170]));
	BUFH_X3M_A12TR DGWClkRightBuff_171(.A(ECK[171]), .Y(DGWClkRightNet[171]));
	BUFH_X3M_A12TR DGWClkRightBuff_172(.A(ECK[172]), .Y(DGWClkRightNet[172]));
	BUFH_X3M_A12TR DGWClkRightBuff_173(.A(ECK[173]), .Y(DGWClkRightNet[173]));
	BUFH_X3M_A12TR DGWClkRightBuff_174(.A(ECK[174]), .Y(DGWClkRightNet[174]));
	BUFH_X3M_A12TR DGWClkRightBuff_175(.A(ECK[175]), .Y(DGWClkRightNet[175]));
	BUFH_X3M_A12TR DGWClkRightBuff_176(.A(ECK[176]), .Y(DGWClkRightNet[176]));
	BUFH_X3M_A12TR DGWClkRightBuff_177(.A(ECK[177]), .Y(DGWClkRightNet[177]));
	BUFH_X3M_A12TR DGWClkRightBuff_178(.A(ECK[178]), .Y(DGWClkRightNet[178]));
	BUFH_X3M_A12TR DGWClkRightBuff_179(.A(ECK[179]), .Y(DGWClkRightNet[179]));
	BUFH_X3M_A12TR DGWClkRightBuff_18(.A(ECK[18]), .Y(DGWClkRightNet[18]));
	BUFH_X3M_A12TR DGWClkRightBuff_180(.A(ECK[180]), .Y(DGWClkRightNet[180]));
	BUFH_X3M_A12TR DGWClkRightBuff_181(.A(ECK[181]), .Y(DGWClkRightNet[181]));
	BUFH_X3M_A12TR DGWClkRightBuff_182(.A(ECK[182]), .Y(DGWClkRightNet[182]));
	BUFH_X3M_A12TR DGWClkRightBuff_183(.A(ECK[183]), .Y(DGWClkRightNet[183]));
	BUFH_X3M_A12TR DGWClkRightBuff_184(.A(ECK[184]), .Y(DGWClkRightNet[184]));
	BUFH_X3M_A12TR DGWClkRightBuff_185(.A(ECK[185]), .Y(DGWClkRightNet[185]));
	BUFH_X3M_A12TR DGWClkRightBuff_186(.A(ECK[186]), .Y(DGWClkRightNet[186]));
	BUFH_X3M_A12TR DGWClkRightBuff_187(.A(ECK[187]), .Y(DGWClkRightNet[187]));
	BUFH_X3M_A12TR DGWClkRightBuff_188(.A(ECK[188]), .Y(DGWClkRightNet[188]));
	BUFH_X3M_A12TR DGWClkRightBuff_189(.A(ECK[189]), .Y(DGWClkRightNet[189]));
	BUFH_X3M_A12TR DGWClkRightBuff_19(.A(ECK[19]), .Y(DGWClkRightNet[19]));
	BUFH_X3M_A12TR DGWClkRightBuff_190(.A(ECK[190]), .Y(DGWClkRightNet[190]));
	BUFH_X3M_A12TR DGWClkRightBuff_191(.A(ECK[191]), .Y(DGWClkRightNet[191]));
	BUFH_X3M_A12TR DGWClkRightBuff_192(.A(ECK[192]), .Y(DGWClkRightNet[192]));
	BUFH_X3M_A12TR DGWClkRightBuff_193(.A(ECK[193]), .Y(DGWClkRightNet[193]));
	BUFH_X3M_A12TR DGWClkRightBuff_194(.A(ECK[194]), .Y(DGWClkRightNet[194]));
	BUFH_X3M_A12TR DGWClkRightBuff_195(.A(ECK[195]), .Y(DGWClkRightNet[195]));
	BUFH_X3M_A12TR DGWClkRightBuff_196(.A(ECK[196]), .Y(DGWClkRightNet[196]));
	BUFH_X3M_A12TR DGWClkRightBuff_197(.A(ECK[197]), .Y(DGWClkRightNet[197]));
	BUFH_X3M_A12TR DGWClkRightBuff_198(.A(ECK[198]), .Y(DGWClkRightNet[198]));
	BUFH_X3M_A12TR DGWClkRightBuff_199(.A(ECK[199]), .Y(DGWClkRightNet[199]));
	BUFH_X3M_A12TR DGWClkRightBuff_2(.A(ECK[2]), .Y(DGWClkRightNet[2]));
	BUFH_X3M_A12TR DGWClkRightBuff_20(.A(ECK[20]), .Y(DGWClkRightNet[20]));
	BUFH_X3M_A12TR DGWClkRightBuff_200(.A(ECK[200]), .Y(DGWClkRightNet[200]));
	BUFH_X3M_A12TR DGWClkRightBuff_201(.A(ECK[201]), .Y(DGWClkRightNet[201]));
	BUFH_X3M_A12TR DGWClkRightBuff_202(.A(ECK[202]), .Y(DGWClkRightNet[202]));
	BUFH_X3M_A12TR DGWClkRightBuff_203(.A(ECK[203]), .Y(DGWClkRightNet[203]));
	BUFH_X3M_A12TR DGWClkRightBuff_204(.A(ECK[204]), .Y(DGWClkRightNet[204]));
	BUFH_X3M_A12TR DGWClkRightBuff_205(.A(ECK[205]), .Y(DGWClkRightNet[205]));
	BUFH_X3M_A12TR DGWClkRightBuff_206(.A(ECK[206]), .Y(DGWClkRightNet[206]));
	BUFH_X3M_A12TR DGWClkRightBuff_207(.A(ECK[207]), .Y(DGWClkRightNet[207]));
	BUFH_X3M_A12TR DGWClkRightBuff_208(.A(ECK[208]), .Y(DGWClkRightNet[208]));
	BUFH_X3M_A12TR DGWClkRightBuff_209(.A(ECK[209]), .Y(DGWClkRightNet[209]));
	BUFH_X3M_A12TR DGWClkRightBuff_21(.A(ECK[21]), .Y(DGWClkRightNet[21]));
	BUFH_X3M_A12TR DGWClkRightBuff_210(.A(ECK[210]), .Y(DGWClkRightNet[210]));
	BUFH_X3M_A12TR DGWClkRightBuff_211(.A(ECK[211]), .Y(DGWClkRightNet[211]));
	BUFH_X3M_A12TR DGWClkRightBuff_212(.A(ECK[212]), .Y(DGWClkRightNet[212]));
	BUFH_X3M_A12TR DGWClkRightBuff_213(.A(ECK[213]), .Y(DGWClkRightNet[213]));
	BUFH_X3M_A12TR DGWClkRightBuff_214(.A(ECK[214]), .Y(DGWClkRightNet[214]));
	BUFH_X3M_A12TR DGWClkRightBuff_215(.A(ECK[215]), .Y(DGWClkRightNet[215]));
	BUFH_X3M_A12TR DGWClkRightBuff_216(.A(ECK[216]), .Y(DGWClkRightNet[216]));
	BUFH_X3M_A12TR DGWClkRightBuff_217(.A(ECK[217]), .Y(DGWClkRightNet[217]));
	BUFH_X3M_A12TR DGWClkRightBuff_218(.A(ECK[218]), .Y(DGWClkRightNet[218]));
	BUFH_X3M_A12TR DGWClkRightBuff_219(.A(ECK[219]), .Y(DGWClkRightNet[219]));
	BUFH_X3M_A12TR DGWClkRightBuff_22(.A(ECK[22]), .Y(DGWClkRightNet[22]));
	BUFH_X3M_A12TR DGWClkRightBuff_220(.A(ECK[220]), .Y(DGWClkRightNet[220]));
	BUFH_X3M_A12TR DGWClkRightBuff_221(.A(ECK[221]), .Y(DGWClkRightNet[221]));
	BUFH_X3M_A12TR DGWClkRightBuff_222(.A(ECK[222]), .Y(DGWClkRightNet[222]));
	BUFH_X3M_A12TR DGWClkRightBuff_223(.A(ECK[223]), .Y(DGWClkRightNet[223]));
	BUFH_X3M_A12TR DGWClkRightBuff_224(.A(ECK[224]), .Y(DGWClkRightNet[224]));
	BUFH_X3M_A12TR DGWClkRightBuff_225(.A(ECK[225]), .Y(DGWClkRightNet[225]));
	BUFH_X3M_A12TR DGWClkRightBuff_226(.A(ECK[226]), .Y(DGWClkRightNet[226]));
	BUFH_X3M_A12TR DGWClkRightBuff_227(.A(ECK[227]), .Y(DGWClkRightNet[227]));
	BUFH_X3M_A12TR DGWClkRightBuff_228(.A(ECK[228]), .Y(DGWClkRightNet[228]));
	BUFH_X3M_A12TR DGWClkRightBuff_229(.A(ECK[229]), .Y(DGWClkRightNet[229]));
	BUFH_X3M_A12TR DGWClkRightBuff_23(.A(ECK[23]), .Y(DGWClkRightNet[23]));
	BUFH_X3M_A12TR DGWClkRightBuff_230(.A(ECK[230]), .Y(DGWClkRightNet[230]));
	BUFH_X3M_A12TR DGWClkRightBuff_231(.A(ECK[231]), .Y(DGWClkRightNet[231]));
	BUFH_X3M_A12TR DGWClkRightBuff_232(.A(ECK[232]), .Y(DGWClkRightNet[232]));
	BUFH_X3M_A12TR DGWClkRightBuff_233(.A(ECK[233]), .Y(DGWClkRightNet[233]));
	BUFH_X3M_A12TR DGWClkRightBuff_234(.A(ECK[234]), .Y(DGWClkRightNet[234]));
	BUFH_X3M_A12TR DGWClkRightBuff_235(.A(ECK[235]), .Y(DGWClkRightNet[235]));
	BUFH_X3M_A12TR DGWClkRightBuff_236(.A(ECK[236]), .Y(DGWClkRightNet[236]));
	BUFH_X3M_A12TR DGWClkRightBuff_237(.A(ECK[237]), .Y(DGWClkRightNet[237]));
	BUFH_X3M_A12TR DGWClkRightBuff_238(.A(ECK[238]), .Y(DGWClkRightNet[238]));
	BUFH_X3M_A12TR DGWClkRightBuff_239(.A(ECK[239]), .Y(DGWClkRightNet[239]));
	BUFH_X3M_A12TR DGWClkRightBuff_24(.A(ECK[24]), .Y(DGWClkRightNet[24]));
	BUFH_X3M_A12TR DGWClkRightBuff_240(.A(ECK[240]), .Y(DGWClkRightNet[240]));
	BUFH_X3M_A12TR DGWClkRightBuff_241(.A(ECK[241]), .Y(DGWClkRightNet[241]));
	BUFH_X3M_A12TR DGWClkRightBuff_242(.A(ECK[242]), .Y(DGWClkRightNet[242]));
	BUFH_X3M_A12TR DGWClkRightBuff_243(.A(ECK[243]), .Y(DGWClkRightNet[243]));
	BUFH_X3M_A12TR DGWClkRightBuff_244(.A(ECK[244]), .Y(DGWClkRightNet[244]));
	BUFH_X3M_A12TR DGWClkRightBuff_245(.A(ECK[245]), .Y(DGWClkRightNet[245]));
	BUFH_X3M_A12TR DGWClkRightBuff_246(.A(ECK[246]), .Y(DGWClkRightNet[246]));
	BUFH_X3M_A12TR DGWClkRightBuff_247(.A(ECK[247]), .Y(DGWClkRightNet[247]));
	BUFH_X3M_A12TR DGWClkRightBuff_248(.A(ECK[248]), .Y(DGWClkRightNet[248]));
	BUFH_X3M_A12TR DGWClkRightBuff_249(.A(ECK[249]), .Y(DGWClkRightNet[249]));
	BUFH_X3M_A12TR DGWClkRightBuff_25(.A(ECK[25]), .Y(DGWClkRightNet[25]));
	BUFH_X3M_A12TR DGWClkRightBuff_250(.A(ECK[250]), .Y(DGWClkRightNet[250]));
	BUFH_X3M_A12TR DGWClkRightBuff_251(.A(ECK[251]), .Y(DGWClkRightNet[251]));
	BUFH_X3M_A12TR DGWClkRightBuff_252(.A(ECK[252]), .Y(DGWClkRightNet[252]));
	BUFH_X3M_A12TR DGWClkRightBuff_253(.A(ECK[253]), .Y(DGWClkRightNet[253]));
	BUFH_X3M_A12TR DGWClkRightBuff_254(.A(ECK[254]), .Y(DGWClkRightNet[254]));
	BUFH_X3M_A12TR DGWClkRightBuff_255(.A(ECK[255]), .Y(DGWClkRightNet[255]));
	BUFH_X3M_A12TR DGWClkRightBuff_26(.A(ECK[26]), .Y(DGWClkRightNet[26]));
	BUFH_X3M_A12TR DGWClkRightBuff_27(.A(ECK[27]), .Y(DGWClkRightNet[27]));
	BUFH_X3M_A12TR DGWClkRightBuff_28(.A(ECK[28]), .Y(DGWClkRightNet[28]));
	BUFH_X3M_A12TR DGWClkRightBuff_29(.A(ECK[29]), .Y(DGWClkRightNet[29]));
	BUFH_X3M_A12TR DGWClkRightBuff_3(.A(ECK[3]), .Y(DGWClkRightNet[3]));
	BUFH_X3M_A12TR DGWClkRightBuff_30(.A(ECK[30]), .Y(DGWClkRightNet[30]));
	BUFH_X3M_A12TR DGWClkRightBuff_31(.A(ECK[31]), .Y(DGWClkRightNet[31]));
	BUFH_X3M_A12TR DGWClkRightBuff_32(.A(ECK[32]), .Y(DGWClkRightNet[32]));
	BUFH_X3M_A12TR DGWClkRightBuff_33(.A(ECK[33]), .Y(DGWClkRightNet[33]));
	BUFH_X3M_A12TR DGWClkRightBuff_34(.A(ECK[34]), .Y(DGWClkRightNet[34]));
	BUFH_X3M_A12TR DGWClkRightBuff_35(.A(ECK[35]), .Y(DGWClkRightNet[35]));
	BUFH_X3M_A12TR DGWClkRightBuff_36(.A(ECK[36]), .Y(DGWClkRightNet[36]));
	BUFH_X3M_A12TR DGWClkRightBuff_37(.A(ECK[37]), .Y(DGWClkRightNet[37]));
	BUFH_X3M_A12TR DGWClkRightBuff_38(.A(ECK[38]), .Y(DGWClkRightNet[38]));
	BUFH_X3M_A12TR DGWClkRightBuff_39(.A(ECK[39]), .Y(DGWClkRightNet[39]));
	BUFH_X3M_A12TR DGWClkRightBuff_4(.A(ECK[4]), .Y(DGWClkRightNet[4]));
	BUFH_X3M_A12TR DGWClkRightBuff_40(.A(ECK[40]), .Y(DGWClkRightNet[40]));
	BUFH_X3M_A12TR DGWClkRightBuff_41(.A(ECK[41]), .Y(DGWClkRightNet[41]));
	BUFH_X3M_A12TR DGWClkRightBuff_42(.A(ECK[42]), .Y(DGWClkRightNet[42]));
	BUFH_X3M_A12TR DGWClkRightBuff_43(.A(ECK[43]), .Y(DGWClkRightNet[43]));
	BUFH_X3M_A12TR DGWClkRightBuff_44(.A(ECK[44]), .Y(DGWClkRightNet[44]));
	BUFH_X3M_A12TR DGWClkRightBuff_45(.A(ECK[45]), .Y(DGWClkRightNet[45]));
	BUFH_X3M_A12TR DGWClkRightBuff_46(.A(ECK[46]), .Y(DGWClkRightNet[46]));
	BUFH_X3M_A12TR DGWClkRightBuff_47(.A(ECK[47]), .Y(DGWClkRightNet[47]));
	BUFH_X3M_A12TR DGWClkRightBuff_48(.A(ECK[48]), .Y(DGWClkRightNet[48]));
	BUFH_X3M_A12TR DGWClkRightBuff_49(.A(ECK[49]), .Y(DGWClkRightNet[49]));
	BUFH_X3M_A12TR DGWClkRightBuff_5(.A(ECK[5]), .Y(DGWClkRightNet[5]));
	BUFH_X3M_A12TR DGWClkRightBuff_50(.A(ECK[50]), .Y(DGWClkRightNet[50]));
	BUFH_X3M_A12TR DGWClkRightBuff_51(.A(ECK[51]), .Y(DGWClkRightNet[51]));
	BUFH_X3M_A12TR DGWClkRightBuff_52(.A(ECK[52]), .Y(DGWClkRightNet[52]));
	BUFH_X3M_A12TR DGWClkRightBuff_53(.A(ECK[53]), .Y(DGWClkRightNet[53]));
	BUFH_X3M_A12TR DGWClkRightBuff_54(.A(ECK[54]), .Y(DGWClkRightNet[54]));
	BUFH_X3M_A12TR DGWClkRightBuff_55(.A(ECK[55]), .Y(DGWClkRightNet[55]));
	BUFH_X3M_A12TR DGWClkRightBuff_56(.A(ECK[56]), .Y(DGWClkRightNet[56]));
	BUFH_X3M_A12TR DGWClkRightBuff_57(.A(ECK[57]), .Y(DGWClkRightNet[57]));
	BUFH_X3M_A12TR DGWClkRightBuff_58(.A(ECK[58]), .Y(DGWClkRightNet[58]));
	BUFH_X3M_A12TR DGWClkRightBuff_59(.A(ECK[59]), .Y(DGWClkRightNet[59]));
	BUFH_X3M_A12TR DGWClkRightBuff_6(.A(ECK[6]), .Y(DGWClkRightNet[6]));
	BUFH_X3M_A12TR DGWClkRightBuff_60(.A(ECK[60]), .Y(DGWClkRightNet[60]));
	BUFH_X3M_A12TR DGWClkRightBuff_61(.A(ECK[61]), .Y(DGWClkRightNet[61]));
	BUFH_X3M_A12TR DGWClkRightBuff_62(.A(ECK[62]), .Y(DGWClkRightNet[62]));
	BUFH_X3M_A12TR DGWClkRightBuff_63(.A(ECK[63]), .Y(DGWClkRightNet[63]));
	BUFH_X3M_A12TR DGWClkRightBuff_64(.A(ECK[64]), .Y(DGWClkRightNet[64]));
	BUFH_X3M_A12TR DGWClkRightBuff_65(.A(ECK[65]), .Y(DGWClkRightNet[65]));
	BUFH_X3M_A12TR DGWClkRightBuff_66(.A(ECK[66]), .Y(DGWClkRightNet[66]));
	BUFH_X3M_A12TR DGWClkRightBuff_67(.A(ECK[67]), .Y(DGWClkRightNet[67]));
	BUFH_X3M_A12TR DGWClkRightBuff_68(.A(ECK[68]), .Y(DGWClkRightNet[68]));
	BUFH_X3M_A12TR DGWClkRightBuff_69(.A(ECK[69]), .Y(DGWClkRightNet[69]));
	BUFH_X3M_A12TR DGWClkRightBuff_7(.A(ECK[7]), .Y(DGWClkRightNet[7]));
	BUFH_X3M_A12TR DGWClkRightBuff_70(.A(ECK[70]), .Y(DGWClkRightNet[70]));
	BUFH_X3M_A12TR DGWClkRightBuff_71(.A(ECK[71]), .Y(DGWClkRightNet[71]));
	BUFH_X3M_A12TR DGWClkRightBuff_72(.A(ECK[72]), .Y(DGWClkRightNet[72]));
	BUFH_X3M_A12TR DGWClkRightBuff_73(.A(ECK[73]), .Y(DGWClkRightNet[73]));
	BUFH_X3M_A12TR DGWClkRightBuff_74(.A(ECK[74]), .Y(DGWClkRightNet[74]));
	BUFH_X3M_A12TR DGWClkRightBuff_75(.A(ECK[75]), .Y(DGWClkRightNet[75]));
	BUFH_X3M_A12TR DGWClkRightBuff_76(.A(ECK[76]), .Y(DGWClkRightNet[76]));
	BUFH_X3M_A12TR DGWClkRightBuff_77(.A(ECK[77]), .Y(DGWClkRightNet[77]));
	BUFH_X3M_A12TR DGWClkRightBuff_78(.A(ECK[78]), .Y(DGWClkRightNet[78]));
	BUFH_X3M_A12TR DGWClkRightBuff_79(.A(ECK[79]), .Y(DGWClkRightNet[79]));
	BUFH_X3M_A12TR DGWClkRightBuff_8(.A(ECK[8]), .Y(DGWClkRightNet[8]));
	BUFH_X3M_A12TR DGWClkRightBuff_80(.A(ECK[80]), .Y(DGWClkRightNet[80]));
	BUFH_X3M_A12TR DGWClkRightBuff_81(.A(ECK[81]), .Y(DGWClkRightNet[81]));
	BUFH_X3M_A12TR DGWClkRightBuff_82(.A(ECK[82]), .Y(DGWClkRightNet[82]));
	BUFH_X3M_A12TR DGWClkRightBuff_83(.A(ECK[83]), .Y(DGWClkRightNet[83]));
	BUFH_X3M_A12TR DGWClkRightBuff_84(.A(ECK[84]), .Y(DGWClkRightNet[84]));
	BUFH_X3M_A12TR DGWClkRightBuff_85(.A(ECK[85]), .Y(DGWClkRightNet[85]));
	BUFH_X3M_A12TR DGWClkRightBuff_86(.A(ECK[86]), .Y(DGWClkRightNet[86]));
	BUFH_X3M_A12TR DGWClkRightBuff_87(.A(ECK[87]), .Y(DGWClkRightNet[87]));
	BUFH_X3M_A12TR DGWClkRightBuff_88(.A(ECK[88]), .Y(DGWClkRightNet[88]));
	BUFH_X3M_A12TR DGWClkRightBuff_89(.A(ECK[89]), .Y(DGWClkRightNet[89]));
	BUFH_X3M_A12TR DGWClkRightBuff_9(.A(ECK[9]), .Y(DGWClkRightNet[9]));
	BUFH_X3M_A12TR DGWClkRightBuff_90(.A(ECK[90]), .Y(DGWClkRightNet[90]));
	BUFH_X3M_A12TR DGWClkRightBuff_91(.A(ECK[91]), .Y(DGWClkRightNet[91]));
	BUFH_X3M_A12TR DGWClkRightBuff_92(.A(ECK[92]), .Y(DGWClkRightNet[92]));
	BUFH_X3M_A12TR DGWClkRightBuff_93(.A(ECK[93]), .Y(DGWClkRightNet[93]));
	BUFH_X3M_A12TR DGWClkRightBuff_94(.A(ECK[94]), .Y(DGWClkRightNet[94]));
	BUFH_X3M_A12TR DGWClkRightBuff_95(.A(ECK[95]), .Y(DGWClkRightNet[95]));
	BUFH_X3M_A12TR DGWClkRightBuff_96(.A(ECK[96]), .Y(DGWClkRightNet[96]));
	BUFH_X3M_A12TR DGWClkRightBuff_97(.A(ECK[97]), .Y(DGWClkRightNet[97]));
	BUFH_X3M_A12TR DGWClkRightBuff_98(.A(ECK[98]), .Y(DGWClkRightNet[98]));
	BUFH_X3M_A12TR DGWClkRightBuff_99(.A(ECK[99]), .Y(DGWClkRightNet[99]));

endmodule
