

module row_decoder (decoder_in, decoder_out);

	//ports
	output [255:0] decoder_out;
	input [7:0] decoder_in;

	//wires
	wire [255:0] decoder_out;
	wire [7:0] decoder_in;
	wire [31:0] PreDec_out;

	//instances
	NOR2_X1A_A12TR PostDec_00(.A(PreDec_out[0]), .B(PreDec_out[16]), .Y(decoder_out[0]));
	NOR2_X1A_A12TR PostDec_01(.A(PreDec_out[1]), .B(PreDec_out[16]), .Y(decoder_out[1]));
	NOR2_X1A_A12TR PostDec_02(.A(PreDec_out[2]), .B(PreDec_out[16]), .Y(decoder_out[2]));
	NOR2_X1A_A12TR PostDec_03(.A(PreDec_out[3]), .B(PreDec_out[16]), .Y(decoder_out[3]));
	NOR2_X1A_A12TR PostDec_04(.A(PreDec_out[4]), .B(PreDec_out[16]), .Y(decoder_out[4]));
	NOR2_X1A_A12TR PostDec_05(.A(PreDec_out[5]), .B(PreDec_out[16]), .Y(decoder_out[5]));
	NOR2_X1A_A12TR PostDec_06(.A(PreDec_out[6]), .B(PreDec_out[16]), .Y(decoder_out[6]));
	NOR2_X1A_A12TR PostDec_07(.A(PreDec_out[7]), .B(PreDec_out[16]), .Y(decoder_out[7]));
	NOR2_X1A_A12TR PostDec_08(.A(PreDec_out[8]), .B(PreDec_out[16]), .Y(decoder_out[8]));
	NOR2_X1A_A12TR PostDec_09(.A(PreDec_out[9]), .B(PreDec_out[16]), .Y(decoder_out[9]));
	NOR2_X1A_A12TR PostDec_10(.A(PreDec_out[10]), .B(PreDec_out[16]), .Y(decoder_out[10]));
	NOR2_X1A_A12TR PostDec_100(.A(PreDec_out[4]), .B(PreDec_out[22]), .Y(decoder_out[100]));
	NOR2_X1A_A12TR PostDec_101(.A(PreDec_out[5]), .B(PreDec_out[22]), .Y(decoder_out[101]));
	NOR2_X1A_A12TR PostDec_102(.A(PreDec_out[6]), .B(PreDec_out[22]), .Y(decoder_out[102]));
	NOR2_X1A_A12TR PostDec_103(.A(PreDec_out[7]), .B(PreDec_out[22]), .Y(decoder_out[103]));
	NOR2_X1A_A12TR PostDec_104(.A(PreDec_out[8]), .B(PreDec_out[22]), .Y(decoder_out[104]));
	NOR2_X1A_A12TR PostDec_105(.A(PreDec_out[9]), .B(PreDec_out[22]), .Y(decoder_out[105]));
	NOR2_X1A_A12TR PostDec_106(.A(PreDec_out[10]), .B(PreDec_out[22]), .Y(decoder_out[106]));
	NOR2_X1A_A12TR PostDec_107(.A(PreDec_out[11]), .B(PreDec_out[22]), .Y(decoder_out[107]));
	NOR2_X1A_A12TR PostDec_108(.A(PreDec_out[12]), .B(PreDec_out[22]), .Y(decoder_out[108]));
	NOR2_X1A_A12TR PostDec_109(.A(PreDec_out[13]), .B(PreDec_out[22]), .Y(decoder_out[109]));
	NOR2_X1A_A12TR PostDec_11(.A(PreDec_out[11]), .B(PreDec_out[16]), .Y(decoder_out[11]));
	NOR2_X1A_A12TR PostDec_110(.A(PreDec_out[14]), .B(PreDec_out[22]), .Y(decoder_out[110]));
	NOR2_X1A_A12TR PostDec_111(.A(PreDec_out[15]), .B(PreDec_out[22]), .Y(decoder_out[111]));
	NOR2_X1A_A12TR PostDec_112(.A(PreDec_out[0]), .B(PreDec_out[23]), .Y(decoder_out[112]));
	NOR2_X1A_A12TR PostDec_113(.A(PreDec_out[1]), .B(PreDec_out[23]), .Y(decoder_out[113]));
	NOR2_X1A_A12TR PostDec_114(.A(PreDec_out[2]), .B(PreDec_out[23]), .Y(decoder_out[114]));
	NOR2_X1A_A12TR PostDec_115(.A(PreDec_out[3]), .B(PreDec_out[23]), .Y(decoder_out[115]));
	NOR2_X1A_A12TR PostDec_116(.A(PreDec_out[4]), .B(PreDec_out[23]), .Y(decoder_out[116]));
	NOR2_X1A_A12TR PostDec_117(.A(PreDec_out[5]), .B(PreDec_out[23]), .Y(decoder_out[117]));
	NOR2_X1A_A12TR PostDec_118(.A(PreDec_out[6]), .B(PreDec_out[23]), .Y(decoder_out[118]));
	NOR2_X1A_A12TR PostDec_119(.A(PreDec_out[7]), .B(PreDec_out[23]), .Y(decoder_out[119]));
	NOR2_X1A_A12TR PostDec_12(.A(PreDec_out[12]), .B(PreDec_out[16]), .Y(decoder_out[12]));
	NOR2_X1A_A12TR PostDec_120(.A(PreDec_out[8]), .B(PreDec_out[23]), .Y(decoder_out[120]));
	NOR2_X1A_A12TR PostDec_121(.A(PreDec_out[9]), .B(PreDec_out[23]), .Y(decoder_out[121]));
	NOR2_X1A_A12TR PostDec_122(.A(PreDec_out[10]), .B(PreDec_out[23]), .Y(decoder_out[122]));
	NOR2_X1A_A12TR PostDec_123(.A(PreDec_out[11]), .B(PreDec_out[23]), .Y(decoder_out[123]));
	NOR2_X1A_A12TR PostDec_124(.A(PreDec_out[12]), .B(PreDec_out[23]), .Y(decoder_out[124]));
	NOR2_X1A_A12TR PostDec_125(.A(PreDec_out[13]), .B(PreDec_out[23]), .Y(decoder_out[125]));
	NOR2_X1A_A12TR PostDec_126(.A(PreDec_out[14]), .B(PreDec_out[23]), .Y(decoder_out[126]));
	NOR2_X1A_A12TR PostDec_127(.A(PreDec_out[15]), .B(PreDec_out[23]), .Y(decoder_out[127]));
	NOR2_X1A_A12TR PostDec_128(.A(PreDec_out[0]), .B(PreDec_out[24]), .Y(decoder_out[128]));
	NOR2_X1A_A12TR PostDec_129(.A(PreDec_out[1]), .B(PreDec_out[24]), .Y(decoder_out[129]));
	NOR2_X1A_A12TR PostDec_13(.A(PreDec_out[13]), .B(PreDec_out[16]), .Y(decoder_out[13]));
	NOR2_X1A_A12TR PostDec_130(.A(PreDec_out[2]), .B(PreDec_out[24]), .Y(decoder_out[130]));
	NOR2_X1A_A12TR PostDec_131(.A(PreDec_out[3]), .B(PreDec_out[24]), .Y(decoder_out[131]));
	NOR2_X1A_A12TR PostDec_132(.A(PreDec_out[4]), .B(PreDec_out[24]), .Y(decoder_out[132]));
	NOR2_X1A_A12TR PostDec_133(.A(PreDec_out[5]), .B(PreDec_out[24]), .Y(decoder_out[133]));
	NOR2_X1A_A12TR PostDec_134(.A(PreDec_out[6]), .B(PreDec_out[24]), .Y(decoder_out[134]));
	NOR2_X1A_A12TR PostDec_135(.A(PreDec_out[7]), .B(PreDec_out[24]), .Y(decoder_out[135]));
	NOR2_X1A_A12TR PostDec_136(.A(PreDec_out[8]), .B(PreDec_out[24]), .Y(decoder_out[136]));
	NOR2_X1A_A12TR PostDec_137(.A(PreDec_out[9]), .B(PreDec_out[24]), .Y(decoder_out[137]));
	NOR2_X1A_A12TR PostDec_138(.A(PreDec_out[10]), .B(PreDec_out[24]), .Y(decoder_out[138]));
	NOR2_X1A_A12TR PostDec_139(.A(PreDec_out[11]), .B(PreDec_out[24]), .Y(decoder_out[139]));
	NOR2_X1A_A12TR PostDec_14(.A(PreDec_out[14]), .B(PreDec_out[16]), .Y(decoder_out[14]));
	NOR2_X1A_A12TR PostDec_140(.A(PreDec_out[12]), .B(PreDec_out[24]), .Y(decoder_out[140]));
	NOR2_X1A_A12TR PostDec_141(.A(PreDec_out[13]), .B(PreDec_out[24]), .Y(decoder_out[141]));
	NOR2_X1A_A12TR PostDec_142(.A(PreDec_out[14]), .B(PreDec_out[24]), .Y(decoder_out[142]));
	NOR2_X1A_A12TR PostDec_143(.A(PreDec_out[15]), .B(PreDec_out[24]), .Y(decoder_out[143]));
	NOR2_X1A_A12TR PostDec_144(.A(PreDec_out[0]), .B(PreDec_out[25]), .Y(decoder_out[144]));
	NOR2_X1A_A12TR PostDec_145(.A(PreDec_out[1]), .B(PreDec_out[25]), .Y(decoder_out[145]));
	NOR2_X1A_A12TR PostDec_146(.A(PreDec_out[2]), .B(PreDec_out[25]), .Y(decoder_out[146]));
	NOR2_X1A_A12TR PostDec_147(.A(PreDec_out[3]), .B(PreDec_out[25]), .Y(decoder_out[147]));
	NOR2_X1A_A12TR PostDec_148(.A(PreDec_out[4]), .B(PreDec_out[25]), .Y(decoder_out[148]));
	NOR2_X1A_A12TR PostDec_149(.A(PreDec_out[5]), .B(PreDec_out[25]), .Y(decoder_out[149]));
	NOR2_X1A_A12TR PostDec_15(.A(PreDec_out[15]), .B(PreDec_out[16]), .Y(decoder_out[15]));
	NOR2_X1A_A12TR PostDec_150(.A(PreDec_out[6]), .B(PreDec_out[25]), .Y(decoder_out[150]));
	NOR2_X1A_A12TR PostDec_151(.A(PreDec_out[7]), .B(PreDec_out[25]), .Y(decoder_out[151]));
	NOR2_X1A_A12TR PostDec_152(.A(PreDec_out[8]), .B(PreDec_out[25]), .Y(decoder_out[152]));
	NOR2_X1A_A12TR PostDec_153(.A(PreDec_out[9]), .B(PreDec_out[25]), .Y(decoder_out[153]));
	NOR2_X1A_A12TR PostDec_154(.A(PreDec_out[10]), .B(PreDec_out[25]), .Y(decoder_out[154]));
	NOR2_X1A_A12TR PostDec_155(.A(PreDec_out[11]), .B(PreDec_out[25]), .Y(decoder_out[155]));
	NOR2_X1A_A12TR PostDec_156(.A(PreDec_out[12]), .B(PreDec_out[25]), .Y(decoder_out[156]));
	NOR2_X1A_A12TR PostDec_157(.A(PreDec_out[13]), .B(PreDec_out[25]), .Y(decoder_out[157]));
	NOR2_X1A_A12TR PostDec_158(.A(PreDec_out[14]), .B(PreDec_out[25]), .Y(decoder_out[158]));
	NOR2_X1A_A12TR PostDec_159(.A(PreDec_out[15]), .B(PreDec_out[25]), .Y(decoder_out[159]));
	NOR2_X1A_A12TR PostDec_16(.A(PreDec_out[0]), .B(PreDec_out[17]), .Y(decoder_out[16]));
	NOR2_X1A_A12TR PostDec_160(.A(PreDec_out[0]), .B(PreDec_out[26]), .Y(decoder_out[160]));
	NOR2_X1A_A12TR PostDec_161(.A(PreDec_out[1]), .B(PreDec_out[26]), .Y(decoder_out[161]));
	NOR2_X1A_A12TR PostDec_162(.A(PreDec_out[2]), .B(PreDec_out[26]), .Y(decoder_out[162]));
	NOR2_X1A_A12TR PostDec_163(.A(PreDec_out[3]), .B(PreDec_out[26]), .Y(decoder_out[163]));
	NOR2_X1A_A12TR PostDec_164(.A(PreDec_out[4]), .B(PreDec_out[26]), .Y(decoder_out[164]));
	NOR2_X1A_A12TR PostDec_165(.A(PreDec_out[5]), .B(PreDec_out[26]), .Y(decoder_out[165]));
	NOR2_X1A_A12TR PostDec_166(.A(PreDec_out[6]), .B(PreDec_out[26]), .Y(decoder_out[166]));
	NOR2_X1A_A12TR PostDec_167(.A(PreDec_out[7]), .B(PreDec_out[26]), .Y(decoder_out[167]));
	NOR2_X1A_A12TR PostDec_168(.A(PreDec_out[8]), .B(PreDec_out[26]), .Y(decoder_out[168]));
	NOR2_X1A_A12TR PostDec_169(.A(PreDec_out[9]), .B(PreDec_out[26]), .Y(decoder_out[169]));
	NOR2_X1A_A12TR PostDec_17(.A(PreDec_out[1]), .B(PreDec_out[17]), .Y(decoder_out[17]));
	NOR2_X1A_A12TR PostDec_170(.A(PreDec_out[10]), .B(PreDec_out[26]), .Y(decoder_out[170]));
	NOR2_X1A_A12TR PostDec_171(.A(PreDec_out[11]), .B(PreDec_out[26]), .Y(decoder_out[171]));
	NOR2_X1A_A12TR PostDec_172(.A(PreDec_out[12]), .B(PreDec_out[26]), .Y(decoder_out[172]));
	NOR2_X1A_A12TR PostDec_173(.A(PreDec_out[13]), .B(PreDec_out[26]), .Y(decoder_out[173]));
	NOR2_X1A_A12TR PostDec_174(.A(PreDec_out[14]), .B(PreDec_out[26]), .Y(decoder_out[174]));
	NOR2_X1A_A12TR PostDec_175(.A(PreDec_out[15]), .B(PreDec_out[26]), .Y(decoder_out[175]));
	NOR2_X1A_A12TR PostDec_176(.A(PreDec_out[0]), .B(PreDec_out[27]), .Y(decoder_out[176]));
	NOR2_X1A_A12TR PostDec_177(.A(PreDec_out[1]), .B(PreDec_out[27]), .Y(decoder_out[177]));
	NOR2_X1A_A12TR PostDec_178(.A(PreDec_out[2]), .B(PreDec_out[27]), .Y(decoder_out[178]));
	NOR2_X1A_A12TR PostDec_179(.A(PreDec_out[3]), .B(PreDec_out[27]), .Y(decoder_out[179]));
	NOR2_X1A_A12TR PostDec_18(.A(PreDec_out[2]), .B(PreDec_out[17]), .Y(decoder_out[18]));
	NOR2_X1A_A12TR PostDec_180(.A(PreDec_out[4]), .B(PreDec_out[27]), .Y(decoder_out[180]));
	NOR2_X1A_A12TR PostDec_181(.A(PreDec_out[5]), .B(PreDec_out[27]), .Y(decoder_out[181]));
	NOR2_X1A_A12TR PostDec_182(.A(PreDec_out[6]), .B(PreDec_out[27]), .Y(decoder_out[182]));
	NOR2_X1A_A12TR PostDec_183(.A(PreDec_out[7]), .B(PreDec_out[27]), .Y(decoder_out[183]));
	NOR2_X1A_A12TR PostDec_184(.A(PreDec_out[8]), .B(PreDec_out[27]), .Y(decoder_out[184]));
	NOR2_X1A_A12TR PostDec_185(.A(PreDec_out[9]), .B(PreDec_out[27]), .Y(decoder_out[185]));
	NOR2_X1A_A12TR PostDec_186(.A(PreDec_out[10]), .B(PreDec_out[27]), .Y(decoder_out[186]));
	NOR2_X1A_A12TR PostDec_187(.A(PreDec_out[11]), .B(PreDec_out[27]), .Y(decoder_out[187]));
	NOR2_X1A_A12TR PostDec_188(.A(PreDec_out[12]), .B(PreDec_out[27]), .Y(decoder_out[188]));
	NOR2_X1A_A12TR PostDec_189(.A(PreDec_out[13]), .B(PreDec_out[27]), .Y(decoder_out[189]));
	NOR2_X1A_A12TR PostDec_19(.A(PreDec_out[3]), .B(PreDec_out[17]), .Y(decoder_out[19]));
	NOR2_X1A_A12TR PostDec_190(.A(PreDec_out[14]), .B(PreDec_out[27]), .Y(decoder_out[190]));
	NOR2_X1A_A12TR PostDec_191(.A(PreDec_out[15]), .B(PreDec_out[27]), .Y(decoder_out[191]));
	NOR2_X1A_A12TR PostDec_192(.A(PreDec_out[0]), .B(PreDec_out[28]), .Y(decoder_out[192]));
	NOR2_X1A_A12TR PostDec_193(.A(PreDec_out[1]), .B(PreDec_out[28]), .Y(decoder_out[193]));
	NOR2_X1A_A12TR PostDec_194(.A(PreDec_out[2]), .B(PreDec_out[28]), .Y(decoder_out[194]));
	NOR2_X1A_A12TR PostDec_195(.A(PreDec_out[3]), .B(PreDec_out[28]), .Y(decoder_out[195]));
	NOR2_X1A_A12TR PostDec_196(.A(PreDec_out[4]), .B(PreDec_out[28]), .Y(decoder_out[196]));
	NOR2_X1A_A12TR PostDec_197(.A(PreDec_out[5]), .B(PreDec_out[28]), .Y(decoder_out[197]));
	NOR2_X1A_A12TR PostDec_198(.A(PreDec_out[6]), .B(PreDec_out[28]), .Y(decoder_out[198]));
	NOR2_X1A_A12TR PostDec_199(.A(PreDec_out[7]), .B(PreDec_out[28]), .Y(decoder_out[199]));
	NOR2_X1A_A12TR PostDec_20(.A(PreDec_out[4]), .B(PreDec_out[17]), .Y(decoder_out[20]));
	NOR2_X1A_A12TR PostDec_200(.A(PreDec_out[8]), .B(PreDec_out[28]), .Y(decoder_out[200]));
	NOR2_X1A_A12TR PostDec_201(.A(PreDec_out[9]), .B(PreDec_out[28]), .Y(decoder_out[201]));
	NOR2_X1A_A12TR PostDec_202(.A(PreDec_out[10]), .B(PreDec_out[28]), .Y(decoder_out[202]));
	NOR2_X1A_A12TR PostDec_203(.A(PreDec_out[11]), .B(PreDec_out[28]), .Y(decoder_out[203]));
	NOR2_X1A_A12TR PostDec_204(.A(PreDec_out[12]), .B(PreDec_out[28]), .Y(decoder_out[204]));
	NOR2_X1A_A12TR PostDec_205(.A(PreDec_out[13]), .B(PreDec_out[28]), .Y(decoder_out[205]));
	NOR2_X1A_A12TR PostDec_206(.A(PreDec_out[14]), .B(PreDec_out[28]), .Y(decoder_out[206]));
	NOR2_X1A_A12TR PostDec_207(.A(PreDec_out[15]), .B(PreDec_out[28]), .Y(decoder_out[207]));
	NOR2_X1A_A12TR PostDec_208(.A(PreDec_out[0]), .B(PreDec_out[29]), .Y(decoder_out[208]));
	NOR2_X1A_A12TR PostDec_209(.A(PreDec_out[1]), .B(PreDec_out[29]), .Y(decoder_out[209]));
	NOR2_X1A_A12TR PostDec_21(.A(PreDec_out[5]), .B(PreDec_out[17]), .Y(decoder_out[21]));
	NOR2_X1A_A12TR PostDec_210(.A(PreDec_out[2]), .B(PreDec_out[29]), .Y(decoder_out[210]));
	NOR2_X1A_A12TR PostDec_211(.A(PreDec_out[3]), .B(PreDec_out[29]), .Y(decoder_out[211]));
	NOR2_X1A_A12TR PostDec_212(.A(PreDec_out[4]), .B(PreDec_out[29]), .Y(decoder_out[212]));
	NOR2_X1A_A12TR PostDec_213(.A(PreDec_out[5]), .B(PreDec_out[29]), .Y(decoder_out[213]));
	NOR2_X1A_A12TR PostDec_214(.A(PreDec_out[6]), .B(PreDec_out[29]), .Y(decoder_out[214]));
	NOR2_X1A_A12TR PostDec_215(.A(PreDec_out[7]), .B(PreDec_out[29]), .Y(decoder_out[215]));
	NOR2_X1A_A12TR PostDec_216(.A(PreDec_out[8]), .B(PreDec_out[29]), .Y(decoder_out[216]));
	NOR2_X1A_A12TR PostDec_217(.A(PreDec_out[9]), .B(PreDec_out[29]), .Y(decoder_out[217]));
	NOR2_X1A_A12TR PostDec_218(.A(PreDec_out[10]), .B(PreDec_out[29]), .Y(decoder_out[218]));
	NOR2_X1A_A12TR PostDec_219(.A(PreDec_out[11]), .B(PreDec_out[29]), .Y(decoder_out[219]));
	NOR2_X1A_A12TR PostDec_22(.A(PreDec_out[6]), .B(PreDec_out[17]), .Y(decoder_out[22]));
	NOR2_X1A_A12TR PostDec_220(.A(PreDec_out[12]), .B(PreDec_out[29]), .Y(decoder_out[220]));
	NOR2_X1A_A12TR PostDec_221(.A(PreDec_out[13]), .B(PreDec_out[29]), .Y(decoder_out[221]));
	NOR2_X1A_A12TR PostDec_222(.A(PreDec_out[14]), .B(PreDec_out[29]), .Y(decoder_out[222]));
	NOR2_X1A_A12TR PostDec_223(.A(PreDec_out[15]), .B(PreDec_out[29]), .Y(decoder_out[223]));
	NOR2_X1A_A12TR PostDec_224(.A(PreDec_out[0]), .B(PreDec_out[30]), .Y(decoder_out[224]));
	NOR2_X1A_A12TR PostDec_225(.A(PreDec_out[1]), .B(PreDec_out[30]), .Y(decoder_out[225]));
	NOR2_X1A_A12TR PostDec_226(.A(PreDec_out[2]), .B(PreDec_out[30]), .Y(decoder_out[226]));
	NOR2_X1A_A12TR PostDec_227(.A(PreDec_out[3]), .B(PreDec_out[30]), .Y(decoder_out[227]));
	NOR2_X1A_A12TR PostDec_228(.A(PreDec_out[4]), .B(PreDec_out[30]), .Y(decoder_out[228]));
	NOR2_X1A_A12TR PostDec_229(.A(PreDec_out[5]), .B(PreDec_out[30]), .Y(decoder_out[229]));
	NOR2_X1A_A12TR PostDec_23(.A(PreDec_out[7]), .B(PreDec_out[17]), .Y(decoder_out[23]));
	NOR2_X1A_A12TR PostDec_230(.A(PreDec_out[6]), .B(PreDec_out[30]), .Y(decoder_out[230]));
	NOR2_X1A_A12TR PostDec_231(.A(PreDec_out[7]), .B(PreDec_out[30]), .Y(decoder_out[231]));
	NOR2_X1A_A12TR PostDec_232(.A(PreDec_out[8]), .B(PreDec_out[30]), .Y(decoder_out[232]));
	NOR2_X1A_A12TR PostDec_233(.A(PreDec_out[9]), .B(PreDec_out[30]), .Y(decoder_out[233]));
	NOR2_X1A_A12TR PostDec_234(.A(PreDec_out[10]), .B(PreDec_out[30]), .Y(decoder_out[234]));
	NOR2_X1A_A12TR PostDec_235(.A(PreDec_out[11]), .B(PreDec_out[30]), .Y(decoder_out[235]));
	NOR2_X1A_A12TR PostDec_236(.A(PreDec_out[12]), .B(PreDec_out[30]), .Y(decoder_out[236]));
	NOR2_X1A_A12TR PostDec_237(.A(PreDec_out[13]), .B(PreDec_out[30]), .Y(decoder_out[237]));
	NOR2_X1A_A12TR PostDec_238(.A(PreDec_out[14]), .B(PreDec_out[30]), .Y(decoder_out[238]));
	NOR2_X1A_A12TR PostDec_239(.A(PreDec_out[15]), .B(PreDec_out[30]), .Y(decoder_out[239]));
	NOR2_X1A_A12TR PostDec_24(.A(PreDec_out[8]), .B(PreDec_out[17]), .Y(decoder_out[24]));
	NOR2_X1A_A12TR PostDec_240(.A(PreDec_out[0]), .B(PreDec_out[31]), .Y(decoder_out[240]));
	NOR2_X1A_A12TR PostDec_241(.A(PreDec_out[1]), .B(PreDec_out[31]), .Y(decoder_out[241]));
	NOR2_X1A_A12TR PostDec_242(.A(PreDec_out[2]), .B(PreDec_out[31]), .Y(decoder_out[242]));
	NOR2_X1A_A12TR PostDec_243(.A(PreDec_out[3]), .B(PreDec_out[31]), .Y(decoder_out[243]));
	NOR2_X1A_A12TR PostDec_244(.A(PreDec_out[4]), .B(PreDec_out[31]), .Y(decoder_out[244]));
	NOR2_X1A_A12TR PostDec_245(.A(PreDec_out[5]), .B(PreDec_out[31]), .Y(decoder_out[245]));
	NOR2_X1A_A12TR PostDec_246(.A(PreDec_out[6]), .B(PreDec_out[31]), .Y(decoder_out[246]));
	NOR2_X1A_A12TR PostDec_247(.A(PreDec_out[7]), .B(PreDec_out[31]), .Y(decoder_out[247]));
	NOR2_X1A_A12TR PostDec_248(.A(PreDec_out[8]), .B(PreDec_out[31]), .Y(decoder_out[248]));
	NOR2_X1A_A12TR PostDec_249(.A(PreDec_out[9]), .B(PreDec_out[31]), .Y(decoder_out[249]));
	NOR2_X1A_A12TR PostDec_25(.A(PreDec_out[9]), .B(PreDec_out[17]), .Y(decoder_out[25]));
	NOR2_X1A_A12TR PostDec_250(.A(PreDec_out[10]), .B(PreDec_out[31]), .Y(decoder_out[250]));
	NOR2_X1A_A12TR PostDec_251(.A(PreDec_out[11]), .B(PreDec_out[31]), .Y(decoder_out[251]));
	NOR2_X1A_A12TR PostDec_252(.A(PreDec_out[12]), .B(PreDec_out[31]), .Y(decoder_out[252]));
	NOR2_X1A_A12TR PostDec_253(.A(PreDec_out[13]), .B(PreDec_out[31]), .Y(decoder_out[253]));
	NOR2_X1A_A12TR PostDec_254(.A(PreDec_out[14]), .B(PreDec_out[31]), .Y(decoder_out[254]));
	NOR2_X1A_A12TR PostDec_255(.A(PreDec_out[15]), .B(PreDec_out[31]), .Y(decoder_out[255]));
	NOR2_X1A_A12TR PostDec_26(.A(PreDec_out[10]), .B(PreDec_out[17]), .Y(decoder_out[26]));
	NOR2_X1A_A12TR PostDec_27(.A(PreDec_out[11]), .B(PreDec_out[17]), .Y(decoder_out[27]));
	NOR2_X1A_A12TR PostDec_28(.A(PreDec_out[12]), .B(PreDec_out[17]), .Y(decoder_out[28]));
	NOR2_X1A_A12TR PostDec_29(.A(PreDec_out[13]), .B(PreDec_out[17]), .Y(decoder_out[29]));
	NOR2_X1A_A12TR PostDec_30(.A(PreDec_out[14]), .B(PreDec_out[17]), .Y(decoder_out[30]));
	NOR2_X1A_A12TR PostDec_31(.A(PreDec_out[15]), .B(PreDec_out[17]), .Y(decoder_out[31]));
	NOR2_X1A_A12TR PostDec_32(.A(PreDec_out[0]), .B(PreDec_out[18]), .Y(decoder_out[32]));
	NOR2_X1A_A12TR PostDec_33(.A(PreDec_out[1]), .B(PreDec_out[18]), .Y(decoder_out[33]));
	NOR2_X1A_A12TR PostDec_34(.A(PreDec_out[2]), .B(PreDec_out[18]), .Y(decoder_out[34]));
	NOR2_X1A_A12TR PostDec_35(.A(PreDec_out[3]), .B(PreDec_out[18]), .Y(decoder_out[35]));
	NOR2_X1A_A12TR PostDec_36(.A(PreDec_out[4]), .B(PreDec_out[18]), .Y(decoder_out[36]));
	NOR2_X1A_A12TR PostDec_37(.A(PreDec_out[5]), .B(PreDec_out[18]), .Y(decoder_out[37]));
	NOR2_X1A_A12TR PostDec_38(.A(PreDec_out[6]), .B(PreDec_out[18]), .Y(decoder_out[38]));
	NOR2_X1A_A12TR PostDec_39(.A(PreDec_out[7]), .B(PreDec_out[18]), .Y(decoder_out[39]));
	NOR2_X1A_A12TR PostDec_40(.A(PreDec_out[8]), .B(PreDec_out[18]), .Y(decoder_out[40]));
	NOR2_X1A_A12TR PostDec_41(.A(PreDec_out[9]), .B(PreDec_out[18]), .Y(decoder_out[41]));
	NOR2_X1A_A12TR PostDec_42(.A(PreDec_out[10]), .B(PreDec_out[18]), .Y(decoder_out[42]));
	NOR2_X1A_A12TR PostDec_43(.A(PreDec_out[11]), .B(PreDec_out[18]), .Y(decoder_out[43]));
	NOR2_X1A_A12TR PostDec_44(.A(PreDec_out[12]), .B(PreDec_out[18]), .Y(decoder_out[44]));
	NOR2_X1A_A12TR PostDec_45(.A(PreDec_out[13]), .B(PreDec_out[18]), .Y(decoder_out[45]));
	NOR2_X1A_A12TR PostDec_46(.A(PreDec_out[14]), .B(PreDec_out[18]), .Y(decoder_out[46]));
	NOR2_X1A_A12TR PostDec_47(.A(PreDec_out[15]), .B(PreDec_out[18]), .Y(decoder_out[47]));
	NOR2_X1A_A12TR PostDec_48(.A(PreDec_out[0]), .B(PreDec_out[19]), .Y(decoder_out[48]));
	NOR2_X1A_A12TR PostDec_49(.A(PreDec_out[1]), .B(PreDec_out[19]), .Y(decoder_out[49]));
	NOR2_X1A_A12TR PostDec_50(.A(PreDec_out[2]), .B(PreDec_out[19]), .Y(decoder_out[50]));
	NOR2_X1A_A12TR PostDec_51(.A(PreDec_out[3]), .B(PreDec_out[19]), .Y(decoder_out[51]));
	NOR2_X1A_A12TR PostDec_52(.A(PreDec_out[4]), .B(PreDec_out[19]), .Y(decoder_out[52]));
	NOR2_X1A_A12TR PostDec_53(.A(PreDec_out[5]), .B(PreDec_out[19]), .Y(decoder_out[53]));
	NOR2_X1A_A12TR PostDec_54(.A(PreDec_out[6]), .B(PreDec_out[19]), .Y(decoder_out[54]));
	NOR2_X1A_A12TR PostDec_55(.A(PreDec_out[7]), .B(PreDec_out[19]), .Y(decoder_out[55]));
	NOR2_X1A_A12TR PostDec_56(.A(PreDec_out[8]), .B(PreDec_out[19]), .Y(decoder_out[56]));
	NOR2_X1A_A12TR PostDec_57(.A(PreDec_out[9]), .B(PreDec_out[19]), .Y(decoder_out[57]));
	NOR2_X1A_A12TR PostDec_58(.A(PreDec_out[10]), .B(PreDec_out[19]), .Y(decoder_out[58]));
	NOR2_X1A_A12TR PostDec_59(.A(PreDec_out[11]), .B(PreDec_out[19]), .Y(decoder_out[59]));
	NOR2_X1A_A12TR PostDec_60(.A(PreDec_out[12]), .B(PreDec_out[19]), .Y(decoder_out[60]));
	NOR2_X1A_A12TR PostDec_61(.A(PreDec_out[13]), .B(PreDec_out[19]), .Y(decoder_out[61]));
	NOR2_X1A_A12TR PostDec_62(.A(PreDec_out[14]), .B(PreDec_out[19]), .Y(decoder_out[62]));
	NOR2_X1A_A12TR PostDec_63(.A(PreDec_out[15]), .B(PreDec_out[19]), .Y(decoder_out[63]));
	NOR2_X1A_A12TR PostDec_64(.A(PreDec_out[0]), .B(PreDec_out[20]), .Y(decoder_out[64]));
	NOR2_X1A_A12TR PostDec_65(.A(PreDec_out[1]), .B(PreDec_out[20]), .Y(decoder_out[65]));
	NOR2_X1A_A12TR PostDec_66(.A(PreDec_out[2]), .B(PreDec_out[20]), .Y(decoder_out[66]));
	NOR2_X1A_A12TR PostDec_67(.A(PreDec_out[3]), .B(PreDec_out[20]), .Y(decoder_out[67]));
	NOR2_X1A_A12TR PostDec_68(.A(PreDec_out[4]), .B(PreDec_out[20]), .Y(decoder_out[68]));
	NOR2_X1A_A12TR PostDec_69(.A(PreDec_out[5]), .B(PreDec_out[20]), .Y(decoder_out[69]));
	NOR2_X1A_A12TR PostDec_70(.A(PreDec_out[6]), .B(PreDec_out[20]), .Y(decoder_out[70]));
	NOR2_X1A_A12TR PostDec_71(.A(PreDec_out[7]), .B(PreDec_out[20]), .Y(decoder_out[71]));
	NOR2_X1A_A12TR PostDec_72(.A(PreDec_out[8]), .B(PreDec_out[20]), .Y(decoder_out[72]));
	NOR2_X1A_A12TR PostDec_73(.A(PreDec_out[9]), .B(PreDec_out[20]), .Y(decoder_out[73]));
	NOR2_X1A_A12TR PostDec_74(.A(PreDec_out[10]), .B(PreDec_out[20]), .Y(decoder_out[74]));
	NOR2_X1A_A12TR PostDec_75(.A(PreDec_out[11]), .B(PreDec_out[20]), .Y(decoder_out[75]));
	NOR2_X1A_A12TR PostDec_76(.A(PreDec_out[12]), .B(PreDec_out[20]), .Y(decoder_out[76]));
	NOR2_X1A_A12TR PostDec_77(.A(PreDec_out[13]), .B(PreDec_out[20]), .Y(decoder_out[77]));
	NOR2_X1A_A12TR PostDec_78(.A(PreDec_out[14]), .B(PreDec_out[20]), .Y(decoder_out[78]));
	NOR2_X1A_A12TR PostDec_79(.A(PreDec_out[15]), .B(PreDec_out[20]), .Y(decoder_out[79]));
	NOR2_X1A_A12TR PostDec_80(.A(PreDec_out[0]), .B(PreDec_out[21]), .Y(decoder_out[80]));
	NOR2_X1A_A12TR PostDec_81(.A(PreDec_out[1]), .B(PreDec_out[21]), .Y(decoder_out[81]));
	NOR2_X1A_A12TR PostDec_82(.A(PreDec_out[2]), .B(PreDec_out[21]), .Y(decoder_out[82]));
	NOR2_X1A_A12TR PostDec_83(.A(PreDec_out[3]), .B(PreDec_out[21]), .Y(decoder_out[83]));
	NOR2_X1A_A12TR PostDec_84(.A(PreDec_out[4]), .B(PreDec_out[21]), .Y(decoder_out[84]));
	NOR2_X1A_A12TR PostDec_85(.A(PreDec_out[5]), .B(PreDec_out[21]), .Y(decoder_out[85]));
	NOR2_X1A_A12TR PostDec_86(.A(PreDec_out[6]), .B(PreDec_out[21]), .Y(decoder_out[86]));
	NOR2_X1A_A12TR PostDec_87(.A(PreDec_out[7]), .B(PreDec_out[21]), .Y(decoder_out[87]));
	NOR2_X1A_A12TR PostDec_88(.A(PreDec_out[8]), .B(PreDec_out[21]), .Y(decoder_out[88]));
	NOR2_X1A_A12TR PostDec_89(.A(PreDec_out[9]), .B(PreDec_out[21]), .Y(decoder_out[89]));
	NOR2_X1A_A12TR PostDec_90(.A(PreDec_out[10]), .B(PreDec_out[21]), .Y(decoder_out[90]));
	NOR2_X1A_A12TR PostDec_91(.A(PreDec_out[11]), .B(PreDec_out[21]), .Y(decoder_out[91]));
	NOR2_X1A_A12TR PostDec_92(.A(PreDec_out[12]), .B(PreDec_out[21]), .Y(decoder_out[92]));
	NOR2_X1A_A12TR PostDec_93(.A(PreDec_out[13]), .B(PreDec_out[21]), .Y(decoder_out[93]));
	NOR2_X1A_A12TR PostDec_94(.A(PreDec_out[14]), .B(PreDec_out[21]), .Y(decoder_out[94]));
	NOR2_X1A_A12TR PostDec_95(.A(PreDec_out[15]), .B(PreDec_out[21]), .Y(decoder_out[95]));
	NOR2_X1A_A12TR PostDec_96(.A(PreDec_out[0]), .B(PreDec_out[22]), .Y(decoder_out[96]));
	NOR2_X1A_A12TR PostDec_97(.A(PreDec_out[1]), .B(PreDec_out[22]), .Y(decoder_out[97]));
	NOR2_X1A_A12TR PostDec_98(.A(PreDec_out[2]), .B(PreDec_out[22]), .Y(decoder_out[98]));
	NOR2_X1A_A12TR PostDec_99(.A(PreDec_out[3]), .B(PreDec_out[22]), .Y(decoder_out[99]));
	PreDecoder_4_16 PreDec_0(.decoder_in({decoder_in[3:0]}), .decoder_out({PreDec_out[15:0]}));
	PreDecoder_4_16 PreDec_1(.decoder_in({decoder_in[7:4]}), .decoder_out({PreDec_out[31:16]}));

endmodule
