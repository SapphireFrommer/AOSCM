

module Decoder_4_16 (decoder_in, decoder_out);

    //ports
    input [3:0] decoder_in;
    output [15:0] decoder_out;

    //wires
    wire [3:0] decoder_in;
    wire [15:0] decoder_out;

    //instances

endmodule
