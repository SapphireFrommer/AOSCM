

module read_mux (DOUT, MemoryLatch, RWL);

	//ports
	input [255:0] MemoryLatch;
	input [255:0] RWL;
	output DOUT;

	//wires
	wire [255:0] RWL;
	wire [255:0] w0;
	wire [31:0] w3;
	wire [7:0] w5;
	wire [0:0] w8;
	wire [63:0] w2;
	wire [15:0] w4;
	wire [255:0] MemoryLatch;
	wire [3:0] w6;
	wire [1:0] w7;
	wire [127:0] w1;
	wire DOUT;

	//instances
	INV_X1B_A12TR inv_out(.A(w8[0]), .Y(DOUT));
	NAND2_X1A_A12TR level_1_0(.A(MemoryLatch[0]), .B(RWL[0]), .Y(w0[0]));
	NAND2_X1A_A12TR level_1_1(.A(MemoryLatch[1]), .B(RWL[1]), .Y(w0[1]));
	NAND2_X1A_A12TR level_1_10(.A(MemoryLatch[10]), .B(RWL[10]), .Y(w0[10]));
	NAND2_X1A_A12TR level_1_100(.A(MemoryLatch[100]), .B(RWL[100]), .Y(w0[100]));
	NAND2_X1A_A12TR level_1_101(.A(MemoryLatch[101]), .B(RWL[101]), .Y(w0[101]));
	NAND2_X1A_A12TR level_1_102(.A(MemoryLatch[102]), .B(RWL[102]), .Y(w0[102]));
	NAND2_X1A_A12TR level_1_103(.A(MemoryLatch[103]), .B(RWL[103]), .Y(w0[103]));
	NAND2_X1A_A12TR level_1_104(.A(MemoryLatch[104]), .B(RWL[104]), .Y(w0[104]));
	NAND2_X1A_A12TR level_1_105(.A(MemoryLatch[105]), .B(RWL[105]), .Y(w0[105]));
	NAND2_X1A_A12TR level_1_106(.A(MemoryLatch[106]), .B(RWL[106]), .Y(w0[106]));
	NAND2_X1A_A12TR level_1_107(.A(MemoryLatch[107]), .B(RWL[107]), .Y(w0[107]));
	NAND2_X1A_A12TR level_1_108(.A(MemoryLatch[108]), .B(RWL[108]), .Y(w0[108]));
	NAND2_X1A_A12TR level_1_109(.A(MemoryLatch[109]), .B(RWL[109]), .Y(w0[109]));
	NAND2_X1A_A12TR level_1_11(.A(MemoryLatch[11]), .B(RWL[11]), .Y(w0[11]));
	NAND2_X1A_A12TR level_1_110(.A(MemoryLatch[110]), .B(RWL[110]), .Y(w0[110]));
	NAND2_X1A_A12TR level_1_111(.A(MemoryLatch[111]), .B(RWL[111]), .Y(w0[111]));
	NAND2_X1A_A12TR level_1_112(.A(MemoryLatch[112]), .B(RWL[112]), .Y(w0[112]));
	NAND2_X1A_A12TR level_1_113(.A(MemoryLatch[113]), .B(RWL[113]), .Y(w0[113]));
	NAND2_X1A_A12TR level_1_114(.A(MemoryLatch[114]), .B(RWL[114]), .Y(w0[114]));
	NAND2_X1A_A12TR level_1_115(.A(MemoryLatch[115]), .B(RWL[115]), .Y(w0[115]));
	NAND2_X1A_A12TR level_1_116(.A(MemoryLatch[116]), .B(RWL[116]), .Y(w0[116]));
	NAND2_X1A_A12TR level_1_117(.A(MemoryLatch[117]), .B(RWL[117]), .Y(w0[117]));
	NAND2_X1A_A12TR level_1_118(.A(MemoryLatch[118]), .B(RWL[118]), .Y(w0[118]));
	NAND2_X1A_A12TR level_1_119(.A(MemoryLatch[119]), .B(RWL[119]), .Y(w0[119]));
	NAND2_X1A_A12TR level_1_12(.A(MemoryLatch[12]), .B(RWL[12]), .Y(w0[12]));
	NAND2_X1A_A12TR level_1_120(.A(MemoryLatch[120]), .B(RWL[120]), .Y(w0[120]));
	NAND2_X1A_A12TR level_1_121(.A(MemoryLatch[121]), .B(RWL[121]), .Y(w0[121]));
	NAND2_X1A_A12TR level_1_122(.A(MemoryLatch[122]), .B(RWL[122]), .Y(w0[122]));
	NAND2_X1A_A12TR level_1_123(.A(MemoryLatch[123]), .B(RWL[123]), .Y(w0[123]));
	NAND2_X1A_A12TR level_1_124(.A(MemoryLatch[124]), .B(RWL[124]), .Y(w0[124]));
	NAND2_X1A_A12TR level_1_125(.A(MemoryLatch[125]), .B(RWL[125]), .Y(w0[125]));
	NAND2_X1A_A12TR level_1_126(.A(MemoryLatch[126]), .B(RWL[126]), .Y(w0[126]));
	NAND2_X1A_A12TR level_1_127(.A(MemoryLatch[127]), .B(RWL[127]), .Y(w0[127]));
	NAND2_X1A_A12TR level_1_128(.A(MemoryLatch[128]), .B(RWL[128]), .Y(w0[128]));
	NAND2_X1A_A12TR level_1_129(.A(MemoryLatch[129]), .B(RWL[129]), .Y(w0[129]));
	NAND2_X1A_A12TR level_1_13(.A(MemoryLatch[13]), .B(RWL[13]), .Y(w0[13]));
	NAND2_X1A_A12TR level_1_130(.A(MemoryLatch[130]), .B(RWL[130]), .Y(w0[130]));
	NAND2_X1A_A12TR level_1_131(.A(MemoryLatch[131]), .B(RWL[131]), .Y(w0[131]));
	NAND2_X1A_A12TR level_1_132(.A(MemoryLatch[132]), .B(RWL[132]), .Y(w0[132]));
	NAND2_X1A_A12TR level_1_133(.A(MemoryLatch[133]), .B(RWL[133]), .Y(w0[133]));
	NAND2_X1A_A12TR level_1_134(.A(MemoryLatch[134]), .B(RWL[134]), .Y(w0[134]));
	NAND2_X1A_A12TR level_1_135(.A(MemoryLatch[135]), .B(RWL[135]), .Y(w0[135]));
	NAND2_X1A_A12TR level_1_136(.A(MemoryLatch[136]), .B(RWL[136]), .Y(w0[136]));
	NAND2_X1A_A12TR level_1_137(.A(MemoryLatch[137]), .B(RWL[137]), .Y(w0[137]));
	NAND2_X1A_A12TR level_1_138(.A(MemoryLatch[138]), .B(RWL[138]), .Y(w0[138]));
	NAND2_X1A_A12TR level_1_139(.A(MemoryLatch[139]), .B(RWL[139]), .Y(w0[139]));
	NAND2_X1A_A12TR level_1_14(.A(MemoryLatch[14]), .B(RWL[14]), .Y(w0[14]));
	NAND2_X1A_A12TR level_1_140(.A(MemoryLatch[140]), .B(RWL[140]), .Y(w0[140]));
	NAND2_X1A_A12TR level_1_141(.A(MemoryLatch[141]), .B(RWL[141]), .Y(w0[141]));
	NAND2_X1A_A12TR level_1_142(.A(MemoryLatch[142]), .B(RWL[142]), .Y(w0[142]));
	NAND2_X1A_A12TR level_1_143(.A(MemoryLatch[143]), .B(RWL[143]), .Y(w0[143]));
	NAND2_X1A_A12TR level_1_144(.A(MemoryLatch[144]), .B(RWL[144]), .Y(w0[144]));
	NAND2_X1A_A12TR level_1_145(.A(MemoryLatch[145]), .B(RWL[145]), .Y(w0[145]));
	NAND2_X1A_A12TR level_1_146(.A(MemoryLatch[146]), .B(RWL[146]), .Y(w0[146]));
	NAND2_X1A_A12TR level_1_147(.A(MemoryLatch[147]), .B(RWL[147]), .Y(w0[147]));
	NAND2_X1A_A12TR level_1_148(.A(MemoryLatch[148]), .B(RWL[148]), .Y(w0[148]));
	NAND2_X1A_A12TR level_1_149(.A(MemoryLatch[149]), .B(RWL[149]), .Y(w0[149]));
	NAND2_X1A_A12TR level_1_15(.A(MemoryLatch[15]), .B(RWL[15]), .Y(w0[15]));
	NAND2_X1A_A12TR level_1_150(.A(MemoryLatch[150]), .B(RWL[150]), .Y(w0[150]));
	NAND2_X1A_A12TR level_1_151(.A(MemoryLatch[151]), .B(RWL[151]), .Y(w0[151]));
	NAND2_X1A_A12TR level_1_152(.A(MemoryLatch[152]), .B(RWL[152]), .Y(w0[152]));
	NAND2_X1A_A12TR level_1_153(.A(MemoryLatch[153]), .B(RWL[153]), .Y(w0[153]));
	NAND2_X1A_A12TR level_1_154(.A(MemoryLatch[154]), .B(RWL[154]), .Y(w0[154]));
	NAND2_X1A_A12TR level_1_155(.A(MemoryLatch[155]), .B(RWL[155]), .Y(w0[155]));
	NAND2_X1A_A12TR level_1_156(.A(MemoryLatch[156]), .B(RWL[156]), .Y(w0[156]));
	NAND2_X1A_A12TR level_1_157(.A(MemoryLatch[157]), .B(RWL[157]), .Y(w0[157]));
	NAND2_X1A_A12TR level_1_158(.A(MemoryLatch[158]), .B(RWL[158]), .Y(w0[158]));
	NAND2_X1A_A12TR level_1_159(.A(MemoryLatch[159]), .B(RWL[159]), .Y(w0[159]));
	NAND2_X1A_A12TR level_1_16(.A(MemoryLatch[16]), .B(RWL[16]), .Y(w0[16]));
	NAND2_X1A_A12TR level_1_160(.A(MemoryLatch[160]), .B(RWL[160]), .Y(w0[160]));
	NAND2_X1A_A12TR level_1_161(.A(MemoryLatch[161]), .B(RWL[161]), .Y(w0[161]));
	NAND2_X1A_A12TR level_1_162(.A(MemoryLatch[162]), .B(RWL[162]), .Y(w0[162]));
	NAND2_X1A_A12TR level_1_163(.A(MemoryLatch[163]), .B(RWL[163]), .Y(w0[163]));
	NAND2_X1A_A12TR level_1_164(.A(MemoryLatch[164]), .B(RWL[164]), .Y(w0[164]));
	NAND2_X1A_A12TR level_1_165(.A(MemoryLatch[165]), .B(RWL[165]), .Y(w0[165]));
	NAND2_X1A_A12TR level_1_166(.A(MemoryLatch[166]), .B(RWL[166]), .Y(w0[166]));
	NAND2_X1A_A12TR level_1_167(.A(MemoryLatch[167]), .B(RWL[167]), .Y(w0[167]));
	NAND2_X1A_A12TR level_1_168(.A(MemoryLatch[168]), .B(RWL[168]), .Y(w0[168]));
	NAND2_X1A_A12TR level_1_169(.A(MemoryLatch[169]), .B(RWL[169]), .Y(w0[169]));
	NAND2_X1A_A12TR level_1_17(.A(MemoryLatch[17]), .B(RWL[17]), .Y(w0[17]));
	NAND2_X1A_A12TR level_1_170(.A(MemoryLatch[170]), .B(RWL[170]), .Y(w0[170]));
	NAND2_X1A_A12TR level_1_171(.A(MemoryLatch[171]), .B(RWL[171]), .Y(w0[171]));
	NAND2_X1A_A12TR level_1_172(.A(MemoryLatch[172]), .B(RWL[172]), .Y(w0[172]));
	NAND2_X1A_A12TR level_1_173(.A(MemoryLatch[173]), .B(RWL[173]), .Y(w0[173]));
	NAND2_X1A_A12TR level_1_174(.A(MemoryLatch[174]), .B(RWL[174]), .Y(w0[174]));
	NAND2_X1A_A12TR level_1_175(.A(MemoryLatch[175]), .B(RWL[175]), .Y(w0[175]));
	NAND2_X1A_A12TR level_1_176(.A(MemoryLatch[176]), .B(RWL[176]), .Y(w0[176]));
	NAND2_X1A_A12TR level_1_177(.A(MemoryLatch[177]), .B(RWL[177]), .Y(w0[177]));
	NAND2_X1A_A12TR level_1_178(.A(MemoryLatch[178]), .B(RWL[178]), .Y(w0[178]));
	NAND2_X1A_A12TR level_1_179(.A(MemoryLatch[179]), .B(RWL[179]), .Y(w0[179]));
	NAND2_X1A_A12TR level_1_18(.A(MemoryLatch[18]), .B(RWL[18]), .Y(w0[18]));
	NAND2_X1A_A12TR level_1_180(.A(MemoryLatch[180]), .B(RWL[180]), .Y(w0[180]));
	NAND2_X1A_A12TR level_1_181(.A(MemoryLatch[181]), .B(RWL[181]), .Y(w0[181]));
	NAND2_X1A_A12TR level_1_182(.A(MemoryLatch[182]), .B(RWL[182]), .Y(w0[182]));
	NAND2_X1A_A12TR level_1_183(.A(MemoryLatch[183]), .B(RWL[183]), .Y(w0[183]));
	NAND2_X1A_A12TR level_1_184(.A(MemoryLatch[184]), .B(RWL[184]), .Y(w0[184]));
	NAND2_X1A_A12TR level_1_185(.A(MemoryLatch[185]), .B(RWL[185]), .Y(w0[185]));
	NAND2_X1A_A12TR level_1_186(.A(MemoryLatch[186]), .B(RWL[186]), .Y(w0[186]));
	NAND2_X1A_A12TR level_1_187(.A(MemoryLatch[187]), .B(RWL[187]), .Y(w0[187]));
	NAND2_X1A_A12TR level_1_188(.A(MemoryLatch[188]), .B(RWL[188]), .Y(w0[188]));
	NAND2_X1A_A12TR level_1_189(.A(MemoryLatch[189]), .B(RWL[189]), .Y(w0[189]));
	NAND2_X1A_A12TR level_1_19(.A(MemoryLatch[19]), .B(RWL[19]), .Y(w0[19]));
	NAND2_X1A_A12TR level_1_190(.A(MemoryLatch[190]), .B(RWL[190]), .Y(w0[190]));
	NAND2_X1A_A12TR level_1_191(.A(MemoryLatch[191]), .B(RWL[191]), .Y(w0[191]));
	NAND2_X1A_A12TR level_1_192(.A(MemoryLatch[192]), .B(RWL[192]), .Y(w0[192]));
	NAND2_X1A_A12TR level_1_193(.A(MemoryLatch[193]), .B(RWL[193]), .Y(w0[193]));
	NAND2_X1A_A12TR level_1_194(.A(MemoryLatch[194]), .B(RWL[194]), .Y(w0[194]));
	NAND2_X1A_A12TR level_1_195(.A(MemoryLatch[195]), .B(RWL[195]), .Y(w0[195]));
	NAND2_X1A_A12TR level_1_196(.A(MemoryLatch[196]), .B(RWL[196]), .Y(w0[196]));
	NAND2_X1A_A12TR level_1_197(.A(MemoryLatch[197]), .B(RWL[197]), .Y(w0[197]));
	NAND2_X1A_A12TR level_1_198(.A(MemoryLatch[198]), .B(RWL[198]), .Y(w0[198]));
	NAND2_X1A_A12TR level_1_199(.A(MemoryLatch[199]), .B(RWL[199]), .Y(w0[199]));
	NAND2_X1A_A12TR level_1_2(.A(MemoryLatch[2]), .B(RWL[2]), .Y(w0[2]));
	NAND2_X1A_A12TR level_1_20(.A(MemoryLatch[20]), .B(RWL[20]), .Y(w0[20]));
	NAND2_X1A_A12TR level_1_200(.A(MemoryLatch[200]), .B(RWL[200]), .Y(w0[200]));
	NAND2_X1A_A12TR level_1_201(.A(MemoryLatch[201]), .B(RWL[201]), .Y(w0[201]));
	NAND2_X1A_A12TR level_1_202(.A(MemoryLatch[202]), .B(RWL[202]), .Y(w0[202]));
	NAND2_X1A_A12TR level_1_203(.A(MemoryLatch[203]), .B(RWL[203]), .Y(w0[203]));
	NAND2_X1A_A12TR level_1_204(.A(MemoryLatch[204]), .B(RWL[204]), .Y(w0[204]));
	NAND2_X1A_A12TR level_1_205(.A(MemoryLatch[205]), .B(RWL[205]), .Y(w0[205]));
	NAND2_X1A_A12TR level_1_206(.A(MemoryLatch[206]), .B(RWL[206]), .Y(w0[206]));
	NAND2_X1A_A12TR level_1_207(.A(MemoryLatch[207]), .B(RWL[207]), .Y(w0[207]));
	NAND2_X1A_A12TR level_1_208(.A(MemoryLatch[208]), .B(RWL[208]), .Y(w0[208]));
	NAND2_X1A_A12TR level_1_209(.A(MemoryLatch[209]), .B(RWL[209]), .Y(w0[209]));
	NAND2_X1A_A12TR level_1_21(.A(MemoryLatch[21]), .B(RWL[21]), .Y(w0[21]));
	NAND2_X1A_A12TR level_1_210(.A(MemoryLatch[210]), .B(RWL[210]), .Y(w0[210]));
	NAND2_X1A_A12TR level_1_211(.A(MemoryLatch[211]), .B(RWL[211]), .Y(w0[211]));
	NAND2_X1A_A12TR level_1_212(.A(MemoryLatch[212]), .B(RWL[212]), .Y(w0[212]));
	NAND2_X1A_A12TR level_1_213(.A(MemoryLatch[213]), .B(RWL[213]), .Y(w0[213]));
	NAND2_X1A_A12TR level_1_214(.A(MemoryLatch[214]), .B(RWL[214]), .Y(w0[214]));
	NAND2_X1A_A12TR level_1_215(.A(MemoryLatch[215]), .B(RWL[215]), .Y(w0[215]));
	NAND2_X1A_A12TR level_1_216(.A(MemoryLatch[216]), .B(RWL[216]), .Y(w0[216]));
	NAND2_X1A_A12TR level_1_217(.A(MemoryLatch[217]), .B(RWL[217]), .Y(w0[217]));
	NAND2_X1A_A12TR level_1_218(.A(MemoryLatch[218]), .B(RWL[218]), .Y(w0[218]));
	NAND2_X1A_A12TR level_1_219(.A(MemoryLatch[219]), .B(RWL[219]), .Y(w0[219]));
	NAND2_X1A_A12TR level_1_22(.A(MemoryLatch[22]), .B(RWL[22]), .Y(w0[22]));
	NAND2_X1A_A12TR level_1_220(.A(MemoryLatch[220]), .B(RWL[220]), .Y(w0[220]));
	NAND2_X1A_A12TR level_1_221(.A(MemoryLatch[221]), .B(RWL[221]), .Y(w0[221]));
	NAND2_X1A_A12TR level_1_222(.A(MemoryLatch[222]), .B(RWL[222]), .Y(w0[222]));
	NAND2_X1A_A12TR level_1_223(.A(MemoryLatch[223]), .B(RWL[223]), .Y(w0[223]));
	NAND2_X1A_A12TR level_1_224(.A(MemoryLatch[224]), .B(RWL[224]), .Y(w0[224]));
	NAND2_X1A_A12TR level_1_225(.A(MemoryLatch[225]), .B(RWL[225]), .Y(w0[225]));
	NAND2_X1A_A12TR level_1_226(.A(MemoryLatch[226]), .B(RWL[226]), .Y(w0[226]));
	NAND2_X1A_A12TR level_1_227(.A(MemoryLatch[227]), .B(RWL[227]), .Y(w0[227]));
	NAND2_X1A_A12TR level_1_228(.A(MemoryLatch[228]), .B(RWL[228]), .Y(w0[228]));
	NAND2_X1A_A12TR level_1_229(.A(MemoryLatch[229]), .B(RWL[229]), .Y(w0[229]));
	NAND2_X1A_A12TR level_1_23(.A(MemoryLatch[23]), .B(RWL[23]), .Y(w0[23]));
	NAND2_X1A_A12TR level_1_230(.A(MemoryLatch[230]), .B(RWL[230]), .Y(w0[230]));
	NAND2_X1A_A12TR level_1_231(.A(MemoryLatch[231]), .B(RWL[231]), .Y(w0[231]));
	NAND2_X1A_A12TR level_1_232(.A(MemoryLatch[232]), .B(RWL[232]), .Y(w0[232]));
	NAND2_X1A_A12TR level_1_233(.A(MemoryLatch[233]), .B(RWL[233]), .Y(w0[233]));
	NAND2_X1A_A12TR level_1_234(.A(MemoryLatch[234]), .B(RWL[234]), .Y(w0[234]));
	NAND2_X1A_A12TR level_1_235(.A(MemoryLatch[235]), .B(RWL[235]), .Y(w0[235]));
	NAND2_X1A_A12TR level_1_236(.A(MemoryLatch[236]), .B(RWL[236]), .Y(w0[236]));
	NAND2_X1A_A12TR level_1_237(.A(MemoryLatch[237]), .B(RWL[237]), .Y(w0[237]));
	NAND2_X1A_A12TR level_1_238(.A(MemoryLatch[238]), .B(RWL[238]), .Y(w0[238]));
	NAND2_X1A_A12TR level_1_239(.A(MemoryLatch[239]), .B(RWL[239]), .Y(w0[239]));
	NAND2_X1A_A12TR level_1_24(.A(MemoryLatch[24]), .B(RWL[24]), .Y(w0[24]));
	NAND2_X1A_A12TR level_1_240(.A(MemoryLatch[240]), .B(RWL[240]), .Y(w0[240]));
	NAND2_X1A_A12TR level_1_241(.A(MemoryLatch[241]), .B(RWL[241]), .Y(w0[241]));
	NAND2_X1A_A12TR level_1_242(.A(MemoryLatch[242]), .B(RWL[242]), .Y(w0[242]));
	NAND2_X1A_A12TR level_1_243(.A(MemoryLatch[243]), .B(RWL[243]), .Y(w0[243]));
	NAND2_X1A_A12TR level_1_244(.A(MemoryLatch[244]), .B(RWL[244]), .Y(w0[244]));
	NAND2_X1A_A12TR level_1_245(.A(MemoryLatch[245]), .B(RWL[245]), .Y(w0[245]));
	NAND2_X1A_A12TR level_1_246(.A(MemoryLatch[246]), .B(RWL[246]), .Y(w0[246]));
	NAND2_X1A_A12TR level_1_247(.A(MemoryLatch[247]), .B(RWL[247]), .Y(w0[247]));
	NAND2_X1A_A12TR level_1_248(.A(MemoryLatch[248]), .B(RWL[248]), .Y(w0[248]));
	NAND2_X1A_A12TR level_1_249(.A(MemoryLatch[249]), .B(RWL[249]), .Y(w0[249]));
	NAND2_X1A_A12TR level_1_25(.A(MemoryLatch[25]), .B(RWL[25]), .Y(w0[25]));
	NAND2_X1A_A12TR level_1_250(.A(MemoryLatch[250]), .B(RWL[250]), .Y(w0[250]));
	NAND2_X1A_A12TR level_1_251(.A(MemoryLatch[251]), .B(RWL[251]), .Y(w0[251]));
	NAND2_X1A_A12TR level_1_252(.A(MemoryLatch[252]), .B(RWL[252]), .Y(w0[252]));
	NAND2_X1A_A12TR level_1_253(.A(MemoryLatch[253]), .B(RWL[253]), .Y(w0[253]));
	NAND2_X1A_A12TR level_1_254(.A(MemoryLatch[254]), .B(RWL[254]), .Y(w0[254]));
	NAND2_X1A_A12TR level_1_255(.A(MemoryLatch[255]), .B(RWL[255]), .Y(w0[255]));
	NAND2_X1A_A12TR level_1_26(.A(MemoryLatch[26]), .B(RWL[26]), .Y(w0[26]));
	NAND2_X1A_A12TR level_1_27(.A(MemoryLatch[27]), .B(RWL[27]), .Y(w0[27]));
	NAND2_X1A_A12TR level_1_28(.A(MemoryLatch[28]), .B(RWL[28]), .Y(w0[28]));
	NAND2_X1A_A12TR level_1_29(.A(MemoryLatch[29]), .B(RWL[29]), .Y(w0[29]));
	NAND2_X1A_A12TR level_1_3(.A(MemoryLatch[3]), .B(RWL[3]), .Y(w0[3]));
	NAND2_X1A_A12TR level_1_30(.A(MemoryLatch[30]), .B(RWL[30]), .Y(w0[30]));
	NAND2_X1A_A12TR level_1_31(.A(MemoryLatch[31]), .B(RWL[31]), .Y(w0[31]));
	NAND2_X1A_A12TR level_1_32(.A(MemoryLatch[32]), .B(RWL[32]), .Y(w0[32]));
	NAND2_X1A_A12TR level_1_33(.A(MemoryLatch[33]), .B(RWL[33]), .Y(w0[33]));
	NAND2_X1A_A12TR level_1_34(.A(MemoryLatch[34]), .B(RWL[34]), .Y(w0[34]));
	NAND2_X1A_A12TR level_1_35(.A(MemoryLatch[35]), .B(RWL[35]), .Y(w0[35]));
	NAND2_X1A_A12TR level_1_36(.A(MemoryLatch[36]), .B(RWL[36]), .Y(w0[36]));
	NAND2_X1A_A12TR level_1_37(.A(MemoryLatch[37]), .B(RWL[37]), .Y(w0[37]));
	NAND2_X1A_A12TR level_1_38(.A(MemoryLatch[38]), .B(RWL[38]), .Y(w0[38]));
	NAND2_X1A_A12TR level_1_39(.A(MemoryLatch[39]), .B(RWL[39]), .Y(w0[39]));
	NAND2_X1A_A12TR level_1_4(.A(MemoryLatch[4]), .B(RWL[4]), .Y(w0[4]));
	NAND2_X1A_A12TR level_1_40(.A(MemoryLatch[40]), .B(RWL[40]), .Y(w0[40]));
	NAND2_X1A_A12TR level_1_41(.A(MemoryLatch[41]), .B(RWL[41]), .Y(w0[41]));
	NAND2_X1A_A12TR level_1_42(.A(MemoryLatch[42]), .B(RWL[42]), .Y(w0[42]));
	NAND2_X1A_A12TR level_1_43(.A(MemoryLatch[43]), .B(RWL[43]), .Y(w0[43]));
	NAND2_X1A_A12TR level_1_44(.A(MemoryLatch[44]), .B(RWL[44]), .Y(w0[44]));
	NAND2_X1A_A12TR level_1_45(.A(MemoryLatch[45]), .B(RWL[45]), .Y(w0[45]));
	NAND2_X1A_A12TR level_1_46(.A(MemoryLatch[46]), .B(RWL[46]), .Y(w0[46]));
	NAND2_X1A_A12TR level_1_47(.A(MemoryLatch[47]), .B(RWL[47]), .Y(w0[47]));
	NAND2_X1A_A12TR level_1_48(.A(MemoryLatch[48]), .B(RWL[48]), .Y(w0[48]));
	NAND2_X1A_A12TR level_1_49(.A(MemoryLatch[49]), .B(RWL[49]), .Y(w0[49]));
	NAND2_X1A_A12TR level_1_5(.A(MemoryLatch[5]), .B(RWL[5]), .Y(w0[5]));
	NAND2_X1A_A12TR level_1_50(.A(MemoryLatch[50]), .B(RWL[50]), .Y(w0[50]));
	NAND2_X1A_A12TR level_1_51(.A(MemoryLatch[51]), .B(RWL[51]), .Y(w0[51]));
	NAND2_X1A_A12TR level_1_52(.A(MemoryLatch[52]), .B(RWL[52]), .Y(w0[52]));
	NAND2_X1A_A12TR level_1_53(.A(MemoryLatch[53]), .B(RWL[53]), .Y(w0[53]));
	NAND2_X1A_A12TR level_1_54(.A(MemoryLatch[54]), .B(RWL[54]), .Y(w0[54]));
	NAND2_X1A_A12TR level_1_55(.A(MemoryLatch[55]), .B(RWL[55]), .Y(w0[55]));
	NAND2_X1A_A12TR level_1_56(.A(MemoryLatch[56]), .B(RWL[56]), .Y(w0[56]));
	NAND2_X1A_A12TR level_1_57(.A(MemoryLatch[57]), .B(RWL[57]), .Y(w0[57]));
	NAND2_X1A_A12TR level_1_58(.A(MemoryLatch[58]), .B(RWL[58]), .Y(w0[58]));
	NAND2_X1A_A12TR level_1_59(.A(MemoryLatch[59]), .B(RWL[59]), .Y(w0[59]));
	NAND2_X1A_A12TR level_1_6(.A(MemoryLatch[6]), .B(RWL[6]), .Y(w0[6]));
	NAND2_X1A_A12TR level_1_60(.A(MemoryLatch[60]), .B(RWL[60]), .Y(w0[60]));
	NAND2_X1A_A12TR level_1_61(.A(MemoryLatch[61]), .B(RWL[61]), .Y(w0[61]));
	NAND2_X1A_A12TR level_1_62(.A(MemoryLatch[62]), .B(RWL[62]), .Y(w0[62]));
	NAND2_X1A_A12TR level_1_63(.A(MemoryLatch[63]), .B(RWL[63]), .Y(w0[63]));
	NAND2_X1A_A12TR level_1_64(.A(MemoryLatch[64]), .B(RWL[64]), .Y(w0[64]));
	NAND2_X1A_A12TR level_1_65(.A(MemoryLatch[65]), .B(RWL[65]), .Y(w0[65]));
	NAND2_X1A_A12TR level_1_66(.A(MemoryLatch[66]), .B(RWL[66]), .Y(w0[66]));
	NAND2_X1A_A12TR level_1_67(.A(MemoryLatch[67]), .B(RWL[67]), .Y(w0[67]));
	NAND2_X1A_A12TR level_1_68(.A(MemoryLatch[68]), .B(RWL[68]), .Y(w0[68]));
	NAND2_X1A_A12TR level_1_69(.A(MemoryLatch[69]), .B(RWL[69]), .Y(w0[69]));
	NAND2_X1A_A12TR level_1_7(.A(MemoryLatch[7]), .B(RWL[7]), .Y(w0[7]));
	NAND2_X1A_A12TR level_1_70(.A(MemoryLatch[70]), .B(RWL[70]), .Y(w0[70]));
	NAND2_X1A_A12TR level_1_71(.A(MemoryLatch[71]), .B(RWL[71]), .Y(w0[71]));
	NAND2_X1A_A12TR level_1_72(.A(MemoryLatch[72]), .B(RWL[72]), .Y(w0[72]));
	NAND2_X1A_A12TR level_1_73(.A(MemoryLatch[73]), .B(RWL[73]), .Y(w0[73]));
	NAND2_X1A_A12TR level_1_74(.A(MemoryLatch[74]), .B(RWL[74]), .Y(w0[74]));
	NAND2_X1A_A12TR level_1_75(.A(MemoryLatch[75]), .B(RWL[75]), .Y(w0[75]));
	NAND2_X1A_A12TR level_1_76(.A(MemoryLatch[76]), .B(RWL[76]), .Y(w0[76]));
	NAND2_X1A_A12TR level_1_77(.A(MemoryLatch[77]), .B(RWL[77]), .Y(w0[77]));
	NAND2_X1A_A12TR level_1_78(.A(MemoryLatch[78]), .B(RWL[78]), .Y(w0[78]));
	NAND2_X1A_A12TR level_1_79(.A(MemoryLatch[79]), .B(RWL[79]), .Y(w0[79]));
	NAND2_X1A_A12TR level_1_8(.A(MemoryLatch[8]), .B(RWL[8]), .Y(w0[8]));
	NAND2_X1A_A12TR level_1_80(.A(MemoryLatch[80]), .B(RWL[80]), .Y(w0[80]));
	NAND2_X1A_A12TR level_1_81(.A(MemoryLatch[81]), .B(RWL[81]), .Y(w0[81]));
	NAND2_X1A_A12TR level_1_82(.A(MemoryLatch[82]), .B(RWL[82]), .Y(w0[82]));
	NAND2_X1A_A12TR level_1_83(.A(MemoryLatch[83]), .B(RWL[83]), .Y(w0[83]));
	NAND2_X1A_A12TR level_1_84(.A(MemoryLatch[84]), .B(RWL[84]), .Y(w0[84]));
	NAND2_X1A_A12TR level_1_85(.A(MemoryLatch[85]), .B(RWL[85]), .Y(w0[85]));
	NAND2_X1A_A12TR level_1_86(.A(MemoryLatch[86]), .B(RWL[86]), .Y(w0[86]));
	NAND2_X1A_A12TR level_1_87(.A(MemoryLatch[87]), .B(RWL[87]), .Y(w0[87]));
	NAND2_X1A_A12TR level_1_88(.A(MemoryLatch[88]), .B(RWL[88]), .Y(w0[88]));
	NAND2_X1A_A12TR level_1_89(.A(MemoryLatch[89]), .B(RWL[89]), .Y(w0[89]));
	NAND2_X1A_A12TR level_1_9(.A(MemoryLatch[9]), .B(RWL[9]), .Y(w0[9]));
	NAND2_X1A_A12TR level_1_90(.A(MemoryLatch[90]), .B(RWL[90]), .Y(w0[90]));
	NAND2_X1A_A12TR level_1_91(.A(MemoryLatch[91]), .B(RWL[91]), .Y(w0[91]));
	NAND2_X1A_A12TR level_1_92(.A(MemoryLatch[92]), .B(RWL[92]), .Y(w0[92]));
	NAND2_X1A_A12TR level_1_93(.A(MemoryLatch[93]), .B(RWL[93]), .Y(w0[93]));
	NAND2_X1A_A12TR level_1_94(.A(MemoryLatch[94]), .B(RWL[94]), .Y(w0[94]));
	NAND2_X1A_A12TR level_1_95(.A(MemoryLatch[95]), .B(RWL[95]), .Y(w0[95]));
	NAND2_X1A_A12TR level_1_96(.A(MemoryLatch[96]), .B(RWL[96]), .Y(w0[96]));
	NAND2_X1A_A12TR level_1_97(.A(MemoryLatch[97]), .B(RWL[97]), .Y(w0[97]));
	NAND2_X1A_A12TR level_1_98(.A(MemoryLatch[98]), .B(RWL[98]), .Y(w0[98]));
	NAND2_X1A_A12TR level_1_99(.A(MemoryLatch[99]), .B(RWL[99]), .Y(w0[99]));
	NAND2_X1A_A12TR level_2_0(.A(w0[0]), .B(w0[1]), .Y(w1[0]));
	NAND2_X1A_A12TR level_2_1(.A(w0[2]), .B(w0[3]), .Y(w1[1]));
	NAND2_X1A_A12TR level_2_10(.A(w0[20]), .B(w0[21]), .Y(w1[10]));
	NAND2_X1A_A12TR level_2_100(.A(w0[200]), .B(w0[201]), .Y(w1[100]));
	NAND2_X1A_A12TR level_2_101(.A(w0[202]), .B(w0[203]), .Y(w1[101]));
	NAND2_X1A_A12TR level_2_102(.A(w0[204]), .B(w0[205]), .Y(w1[102]));
	NAND2_X1A_A12TR level_2_103(.A(w0[206]), .B(w0[207]), .Y(w1[103]));
	NAND2_X1A_A12TR level_2_104(.A(w0[208]), .B(w0[209]), .Y(w1[104]));
	NAND2_X1A_A12TR level_2_105(.A(w0[210]), .B(w0[211]), .Y(w1[105]));
	NAND2_X1A_A12TR level_2_106(.A(w0[212]), .B(w0[213]), .Y(w1[106]));
	NAND2_X1A_A12TR level_2_107(.A(w0[214]), .B(w0[215]), .Y(w1[107]));
	NAND2_X1A_A12TR level_2_108(.A(w0[216]), .B(w0[217]), .Y(w1[108]));
	NAND2_X1A_A12TR level_2_109(.A(w0[218]), .B(w0[219]), .Y(w1[109]));
	NAND2_X1A_A12TR level_2_11(.A(w0[22]), .B(w0[23]), .Y(w1[11]));
	NAND2_X1A_A12TR level_2_110(.A(w0[220]), .B(w0[221]), .Y(w1[110]));
	NAND2_X1A_A12TR level_2_111(.A(w0[222]), .B(w0[223]), .Y(w1[111]));
	NAND2_X1A_A12TR level_2_112(.A(w0[224]), .B(w0[225]), .Y(w1[112]));
	NAND2_X1A_A12TR level_2_113(.A(w0[226]), .B(w0[227]), .Y(w1[113]));
	NAND2_X1A_A12TR level_2_114(.A(w0[228]), .B(w0[229]), .Y(w1[114]));
	NAND2_X1A_A12TR level_2_115(.A(w0[230]), .B(w0[231]), .Y(w1[115]));
	NAND2_X1A_A12TR level_2_116(.A(w0[232]), .B(w0[233]), .Y(w1[116]));
	NAND2_X1A_A12TR level_2_117(.A(w0[234]), .B(w0[235]), .Y(w1[117]));
	NAND2_X1A_A12TR level_2_118(.A(w0[236]), .B(w0[237]), .Y(w1[118]));
	NAND2_X1A_A12TR level_2_119(.A(w0[238]), .B(w0[239]), .Y(w1[119]));
	NAND2_X1A_A12TR level_2_12(.A(w0[24]), .B(w0[25]), .Y(w1[12]));
	NAND2_X1A_A12TR level_2_120(.A(w0[240]), .B(w0[241]), .Y(w1[120]));
	NAND2_X1A_A12TR level_2_121(.A(w0[242]), .B(w0[243]), .Y(w1[121]));
	NAND2_X1A_A12TR level_2_122(.A(w0[244]), .B(w0[245]), .Y(w1[122]));
	NAND2_X1A_A12TR level_2_123(.A(w0[246]), .B(w0[247]), .Y(w1[123]));
	NAND2_X1A_A12TR level_2_124(.A(w0[248]), .B(w0[249]), .Y(w1[124]));
	NAND2_X1A_A12TR level_2_125(.A(w0[250]), .B(w0[251]), .Y(w1[125]));
	NAND2_X1A_A12TR level_2_126(.A(w0[252]), .B(w0[253]), .Y(w1[126]));
	NAND2_X1A_A12TR level_2_127(.A(w0[254]), .B(w0[255]), .Y(w1[127]));
	NAND2_X1A_A12TR level_2_13(.A(w0[26]), .B(w0[27]), .Y(w1[13]));
	NAND2_X1A_A12TR level_2_14(.A(w0[28]), .B(w0[29]), .Y(w1[14]));
	NAND2_X1A_A12TR level_2_15(.A(w0[30]), .B(w0[31]), .Y(w1[15]));
	NAND2_X1A_A12TR level_2_16(.A(w0[32]), .B(w0[33]), .Y(w1[16]));
	NAND2_X1A_A12TR level_2_17(.A(w0[34]), .B(w0[35]), .Y(w1[17]));
	NAND2_X1A_A12TR level_2_18(.A(w0[36]), .B(w0[37]), .Y(w1[18]));
	NAND2_X1A_A12TR level_2_19(.A(w0[38]), .B(w0[39]), .Y(w1[19]));
	NAND2_X1A_A12TR level_2_2(.A(w0[4]), .B(w0[5]), .Y(w1[2]));
	NAND2_X1A_A12TR level_2_20(.A(w0[40]), .B(w0[41]), .Y(w1[20]));
	NAND2_X1A_A12TR level_2_21(.A(w0[42]), .B(w0[43]), .Y(w1[21]));
	NAND2_X1A_A12TR level_2_22(.A(w0[44]), .B(w0[45]), .Y(w1[22]));
	NAND2_X1A_A12TR level_2_23(.A(w0[46]), .B(w0[47]), .Y(w1[23]));
	NAND2_X1A_A12TR level_2_24(.A(w0[48]), .B(w0[49]), .Y(w1[24]));
	NAND2_X1A_A12TR level_2_25(.A(w0[50]), .B(w0[51]), .Y(w1[25]));
	NAND2_X1A_A12TR level_2_26(.A(w0[52]), .B(w0[53]), .Y(w1[26]));
	NAND2_X1A_A12TR level_2_27(.A(w0[54]), .B(w0[55]), .Y(w1[27]));
	NAND2_X1A_A12TR level_2_28(.A(w0[56]), .B(w0[57]), .Y(w1[28]));
	NAND2_X1A_A12TR level_2_29(.A(w0[58]), .B(w0[59]), .Y(w1[29]));
	NAND2_X1A_A12TR level_2_3(.A(w0[6]), .B(w0[7]), .Y(w1[3]));
	NAND2_X1A_A12TR level_2_30(.A(w0[60]), .B(w0[61]), .Y(w1[30]));
	NAND2_X1A_A12TR level_2_31(.A(w0[62]), .B(w0[63]), .Y(w1[31]));
	NAND2_X1A_A12TR level_2_32(.A(w0[64]), .B(w0[65]), .Y(w1[32]));
	NAND2_X1A_A12TR level_2_33(.A(w0[66]), .B(w0[67]), .Y(w1[33]));
	NAND2_X1A_A12TR level_2_34(.A(w0[68]), .B(w0[69]), .Y(w1[34]));
	NAND2_X1A_A12TR level_2_35(.A(w0[70]), .B(w0[71]), .Y(w1[35]));
	NAND2_X1A_A12TR level_2_36(.A(w0[72]), .B(w0[73]), .Y(w1[36]));
	NAND2_X1A_A12TR level_2_37(.A(w0[74]), .B(w0[75]), .Y(w1[37]));
	NAND2_X1A_A12TR level_2_38(.A(w0[76]), .B(w0[77]), .Y(w1[38]));
	NAND2_X1A_A12TR level_2_39(.A(w0[78]), .B(w0[79]), .Y(w1[39]));
	NAND2_X1A_A12TR level_2_4(.A(w0[8]), .B(w0[9]), .Y(w1[4]));
	NAND2_X1A_A12TR level_2_40(.A(w0[80]), .B(w0[81]), .Y(w1[40]));
	NAND2_X1A_A12TR level_2_41(.A(w0[82]), .B(w0[83]), .Y(w1[41]));
	NAND2_X1A_A12TR level_2_42(.A(w0[84]), .B(w0[85]), .Y(w1[42]));
	NAND2_X1A_A12TR level_2_43(.A(w0[86]), .B(w0[87]), .Y(w1[43]));
	NAND2_X1A_A12TR level_2_44(.A(w0[88]), .B(w0[89]), .Y(w1[44]));
	NAND2_X1A_A12TR level_2_45(.A(w0[90]), .B(w0[91]), .Y(w1[45]));
	NAND2_X1A_A12TR level_2_46(.A(w0[92]), .B(w0[93]), .Y(w1[46]));
	NAND2_X1A_A12TR level_2_47(.A(w0[94]), .B(w0[95]), .Y(w1[47]));
	NAND2_X1A_A12TR level_2_48(.A(w0[96]), .B(w0[97]), .Y(w1[48]));
	NAND2_X1A_A12TR level_2_49(.A(w0[98]), .B(w0[99]), .Y(w1[49]));
	NAND2_X1A_A12TR level_2_5(.A(w0[10]), .B(w0[11]), .Y(w1[5]));
	NAND2_X1A_A12TR level_2_50(.A(w0[100]), .B(w0[101]), .Y(w1[50]));
	NAND2_X1A_A12TR level_2_51(.A(w0[102]), .B(w0[103]), .Y(w1[51]));
	NAND2_X1A_A12TR level_2_52(.A(w0[104]), .B(w0[105]), .Y(w1[52]));
	NAND2_X1A_A12TR level_2_53(.A(w0[106]), .B(w0[107]), .Y(w1[53]));
	NAND2_X1A_A12TR level_2_54(.A(w0[108]), .B(w0[109]), .Y(w1[54]));
	NAND2_X1A_A12TR level_2_55(.A(w0[110]), .B(w0[111]), .Y(w1[55]));
	NAND2_X1A_A12TR level_2_56(.A(w0[112]), .B(w0[113]), .Y(w1[56]));
	NAND2_X1A_A12TR level_2_57(.A(w0[114]), .B(w0[115]), .Y(w1[57]));
	NAND2_X1A_A12TR level_2_58(.A(w0[116]), .B(w0[117]), .Y(w1[58]));
	NAND2_X1A_A12TR level_2_59(.A(w0[118]), .B(w0[119]), .Y(w1[59]));
	NAND2_X1A_A12TR level_2_6(.A(w0[12]), .B(w0[13]), .Y(w1[6]));
	NAND2_X1A_A12TR level_2_60(.A(w0[120]), .B(w0[121]), .Y(w1[60]));
	NAND2_X1A_A12TR level_2_61(.A(w0[122]), .B(w0[123]), .Y(w1[61]));
	NAND2_X1A_A12TR level_2_62(.A(w0[124]), .B(w0[125]), .Y(w1[62]));
	NAND2_X1A_A12TR level_2_63(.A(w0[126]), .B(w0[127]), .Y(w1[63]));
	NAND2_X1A_A12TR level_2_64(.A(w0[128]), .B(w0[129]), .Y(w1[64]));
	NAND2_X1A_A12TR level_2_65(.A(w0[130]), .B(w0[131]), .Y(w1[65]));
	NAND2_X1A_A12TR level_2_66(.A(w0[132]), .B(w0[133]), .Y(w1[66]));
	NAND2_X1A_A12TR level_2_67(.A(w0[134]), .B(w0[135]), .Y(w1[67]));
	NAND2_X1A_A12TR level_2_68(.A(w0[136]), .B(w0[137]), .Y(w1[68]));
	NAND2_X1A_A12TR level_2_69(.A(w0[138]), .B(w0[139]), .Y(w1[69]));
	NAND2_X1A_A12TR level_2_7(.A(w0[14]), .B(w0[15]), .Y(w1[7]));
	NAND2_X1A_A12TR level_2_70(.A(w0[140]), .B(w0[141]), .Y(w1[70]));
	NAND2_X1A_A12TR level_2_71(.A(w0[142]), .B(w0[143]), .Y(w1[71]));
	NAND2_X1A_A12TR level_2_72(.A(w0[144]), .B(w0[145]), .Y(w1[72]));
	NAND2_X1A_A12TR level_2_73(.A(w0[146]), .B(w0[147]), .Y(w1[73]));
	NAND2_X1A_A12TR level_2_74(.A(w0[148]), .B(w0[149]), .Y(w1[74]));
	NAND2_X1A_A12TR level_2_75(.A(w0[150]), .B(w0[151]), .Y(w1[75]));
	NAND2_X1A_A12TR level_2_76(.A(w0[152]), .B(w0[153]), .Y(w1[76]));
	NAND2_X1A_A12TR level_2_77(.A(w0[154]), .B(w0[155]), .Y(w1[77]));
	NAND2_X1A_A12TR level_2_78(.A(w0[156]), .B(w0[157]), .Y(w1[78]));
	NAND2_X1A_A12TR level_2_79(.A(w0[158]), .B(w0[159]), .Y(w1[79]));
	NAND2_X1A_A12TR level_2_8(.A(w0[16]), .B(w0[17]), .Y(w1[8]));
	NAND2_X1A_A12TR level_2_80(.A(w0[160]), .B(w0[161]), .Y(w1[80]));
	NAND2_X1A_A12TR level_2_81(.A(w0[162]), .B(w0[163]), .Y(w1[81]));
	NAND2_X1A_A12TR level_2_82(.A(w0[164]), .B(w0[165]), .Y(w1[82]));
	NAND2_X1A_A12TR level_2_83(.A(w0[166]), .B(w0[167]), .Y(w1[83]));
	NAND2_X1A_A12TR level_2_84(.A(w0[168]), .B(w0[169]), .Y(w1[84]));
	NAND2_X1A_A12TR level_2_85(.A(w0[170]), .B(w0[171]), .Y(w1[85]));
	NAND2_X1A_A12TR level_2_86(.A(w0[172]), .B(w0[173]), .Y(w1[86]));
	NAND2_X1A_A12TR level_2_87(.A(w0[174]), .B(w0[175]), .Y(w1[87]));
	NAND2_X1A_A12TR level_2_88(.A(w0[176]), .B(w0[177]), .Y(w1[88]));
	NAND2_X1A_A12TR level_2_89(.A(w0[178]), .B(w0[179]), .Y(w1[89]));
	NAND2_X1A_A12TR level_2_9(.A(w0[18]), .B(w0[19]), .Y(w1[9]));
	NAND2_X1A_A12TR level_2_90(.A(w0[180]), .B(w0[181]), .Y(w1[90]));
	NAND2_X1A_A12TR level_2_91(.A(w0[182]), .B(w0[183]), .Y(w1[91]));
	NAND2_X1A_A12TR level_2_92(.A(w0[184]), .B(w0[185]), .Y(w1[92]));
	NAND2_X1A_A12TR level_2_93(.A(w0[186]), .B(w0[187]), .Y(w1[93]));
	NAND2_X1A_A12TR level_2_94(.A(w0[188]), .B(w0[189]), .Y(w1[94]));
	NAND2_X1A_A12TR level_2_95(.A(w0[190]), .B(w0[191]), .Y(w1[95]));
	NAND2_X1A_A12TR level_2_96(.A(w0[192]), .B(w0[193]), .Y(w1[96]));
	NAND2_X1A_A12TR level_2_97(.A(w0[194]), .B(w0[195]), .Y(w1[97]));
	NAND2_X1A_A12TR level_2_98(.A(w0[196]), .B(w0[197]), .Y(w1[98]));
	NAND2_X1A_A12TR level_2_99(.A(w0[198]), .B(w0[199]), .Y(w1[99]));
	NOR2_X1A_A12TR level_3_0(.A(w1[0]), .B(w1[1]), .Y(w2[0]));
	NOR2_X1A_A12TR level_3_1(.A(w1[2]), .B(w1[3]), .Y(w2[1]));
	NOR2_X1A_A12TR level_3_10(.A(w1[20]), .B(w1[21]), .Y(w2[10]));
	NOR2_X1A_A12TR level_3_11(.A(w1[22]), .B(w1[23]), .Y(w2[11]));
	NOR2_X1A_A12TR level_3_12(.A(w1[24]), .B(w1[25]), .Y(w2[12]));
	NOR2_X1A_A12TR level_3_13(.A(w1[26]), .B(w1[27]), .Y(w2[13]));
	NOR2_X1A_A12TR level_3_14(.A(w1[28]), .B(w1[29]), .Y(w2[14]));
	NOR2_X1A_A12TR level_3_15(.A(w1[30]), .B(w1[31]), .Y(w2[15]));
	NOR2_X1A_A12TR level_3_16(.A(w1[32]), .B(w1[33]), .Y(w2[16]));
	NOR2_X1A_A12TR level_3_17(.A(w1[34]), .B(w1[35]), .Y(w2[17]));
	NOR2_X1A_A12TR level_3_18(.A(w1[36]), .B(w1[37]), .Y(w2[18]));
	NOR2_X1A_A12TR level_3_19(.A(w1[38]), .B(w1[39]), .Y(w2[19]));
	NOR2_X1A_A12TR level_3_2(.A(w1[4]), .B(w1[5]), .Y(w2[2]));
	NOR2_X1A_A12TR level_3_20(.A(w1[40]), .B(w1[41]), .Y(w2[20]));
	NOR2_X1A_A12TR level_3_21(.A(w1[42]), .B(w1[43]), .Y(w2[21]));
	NOR2_X1A_A12TR level_3_22(.A(w1[44]), .B(w1[45]), .Y(w2[22]));
	NOR2_X1A_A12TR level_3_23(.A(w1[46]), .B(w1[47]), .Y(w2[23]));
	NOR2_X1A_A12TR level_3_24(.A(w1[48]), .B(w1[49]), .Y(w2[24]));
	NOR2_X1A_A12TR level_3_25(.A(w1[50]), .B(w1[51]), .Y(w2[25]));
	NOR2_X1A_A12TR level_3_26(.A(w1[52]), .B(w1[53]), .Y(w2[26]));
	NOR2_X1A_A12TR level_3_27(.A(w1[54]), .B(w1[55]), .Y(w2[27]));
	NOR2_X1A_A12TR level_3_28(.A(w1[56]), .B(w1[57]), .Y(w2[28]));
	NOR2_X1A_A12TR level_3_29(.A(w1[58]), .B(w1[59]), .Y(w2[29]));
	NOR2_X1A_A12TR level_3_3(.A(w1[6]), .B(w1[7]), .Y(w2[3]));
	NOR2_X1A_A12TR level_3_30(.A(w1[60]), .B(w1[61]), .Y(w2[30]));
	NOR2_X1A_A12TR level_3_31(.A(w1[62]), .B(w1[63]), .Y(w2[31]));
	NOR2_X1A_A12TR level_3_32(.A(w1[64]), .B(w1[65]), .Y(w2[32]));
	NOR2_X1A_A12TR level_3_33(.A(w1[66]), .B(w1[67]), .Y(w2[33]));
	NOR2_X1A_A12TR level_3_34(.A(w1[68]), .B(w1[69]), .Y(w2[34]));
	NOR2_X1A_A12TR level_3_35(.A(w1[70]), .B(w1[71]), .Y(w2[35]));
	NOR2_X1A_A12TR level_3_36(.A(w1[72]), .B(w1[73]), .Y(w2[36]));
	NOR2_X1A_A12TR level_3_37(.A(w1[74]), .B(w1[75]), .Y(w2[37]));
	NOR2_X1A_A12TR level_3_38(.A(w1[76]), .B(w1[77]), .Y(w2[38]));
	NOR2_X1A_A12TR level_3_39(.A(w1[78]), .B(w1[79]), .Y(w2[39]));
	NOR2_X1A_A12TR level_3_4(.A(w1[8]), .B(w1[9]), .Y(w2[4]));
	NOR2_X1A_A12TR level_3_40(.A(w1[80]), .B(w1[81]), .Y(w2[40]));
	NOR2_X1A_A12TR level_3_41(.A(w1[82]), .B(w1[83]), .Y(w2[41]));
	NOR2_X1A_A12TR level_3_42(.A(w1[84]), .B(w1[85]), .Y(w2[42]));
	NOR2_X1A_A12TR level_3_43(.A(w1[86]), .B(w1[87]), .Y(w2[43]));
	NOR2_X1A_A12TR level_3_44(.A(w1[88]), .B(w1[89]), .Y(w2[44]));
	NOR2_X1A_A12TR level_3_45(.A(w1[90]), .B(w1[91]), .Y(w2[45]));
	NOR2_X1A_A12TR level_3_46(.A(w1[92]), .B(w1[93]), .Y(w2[46]));
	NOR2_X1A_A12TR level_3_47(.A(w1[94]), .B(w1[95]), .Y(w2[47]));
	NOR2_X1A_A12TR level_3_48(.A(w1[96]), .B(w1[97]), .Y(w2[48]));
	NOR2_X1A_A12TR level_3_49(.A(w1[98]), .B(w1[99]), .Y(w2[49]));
	NOR2_X1A_A12TR level_3_5(.A(w1[10]), .B(w1[11]), .Y(w2[5]));
	NOR2_X1A_A12TR level_3_50(.A(w1[100]), .B(w1[101]), .Y(w2[50]));
	NOR2_X1A_A12TR level_3_51(.A(w1[102]), .B(w1[103]), .Y(w2[51]));
	NOR2_X1A_A12TR level_3_52(.A(w1[104]), .B(w1[105]), .Y(w2[52]));
	NOR2_X1A_A12TR level_3_53(.A(w1[106]), .B(w1[107]), .Y(w2[53]));
	NOR2_X1A_A12TR level_3_54(.A(w1[108]), .B(w1[109]), .Y(w2[54]));
	NOR2_X1A_A12TR level_3_55(.A(w1[110]), .B(w1[111]), .Y(w2[55]));
	NOR2_X1A_A12TR level_3_56(.A(w1[112]), .B(w1[113]), .Y(w2[56]));
	NOR2_X1A_A12TR level_3_57(.A(w1[114]), .B(w1[115]), .Y(w2[57]));
	NOR2_X1A_A12TR level_3_58(.A(w1[116]), .B(w1[117]), .Y(w2[58]));
	NOR2_X1A_A12TR level_3_59(.A(w1[118]), .B(w1[119]), .Y(w2[59]));
	NOR2_X1A_A12TR level_3_6(.A(w1[12]), .B(w1[13]), .Y(w2[6]));
	NOR2_X1A_A12TR level_3_60(.A(w1[120]), .B(w1[121]), .Y(w2[60]));
	NOR2_X1A_A12TR level_3_61(.A(w1[122]), .B(w1[123]), .Y(w2[61]));
	NOR2_X1A_A12TR level_3_62(.A(w1[124]), .B(w1[125]), .Y(w2[62]));
	NOR2_X1A_A12TR level_3_63(.A(w1[126]), .B(w1[127]), .Y(w2[63]));
	NOR2_X1A_A12TR level_3_7(.A(w1[14]), .B(w1[15]), .Y(w2[7]));
	NOR2_X1A_A12TR level_3_8(.A(w1[16]), .B(w1[17]), .Y(w2[8]));
	NOR2_X1A_A12TR level_3_9(.A(w1[18]), .B(w1[19]), .Y(w2[9]));
	NAND2_X1A_A12TR level_4_0(.A(w2[0]), .B(w2[1]), .Y(w3[0]));
	NAND2_X1A_A12TR level_4_1(.A(w2[2]), .B(w2[3]), .Y(w3[1]));
	NAND2_X1A_A12TR level_4_10(.A(w2[20]), .B(w2[21]), .Y(w3[10]));
	NAND2_X1A_A12TR level_4_11(.A(w2[22]), .B(w2[23]), .Y(w3[11]));
	NAND2_X1A_A12TR level_4_12(.A(w2[24]), .B(w2[25]), .Y(w3[12]));
	NAND2_X1A_A12TR level_4_13(.A(w2[26]), .B(w2[27]), .Y(w3[13]));
	NAND2_X1A_A12TR level_4_14(.A(w2[28]), .B(w2[29]), .Y(w3[14]));
	NAND2_X1A_A12TR level_4_15(.A(w2[30]), .B(w2[31]), .Y(w3[15]));
	NAND2_X1A_A12TR level_4_16(.A(w2[32]), .B(w2[33]), .Y(w3[16]));
	NAND2_X1A_A12TR level_4_17(.A(w2[34]), .B(w2[35]), .Y(w3[17]));
	NAND2_X1A_A12TR level_4_18(.A(w2[36]), .B(w2[37]), .Y(w3[18]));
	NAND2_X1A_A12TR level_4_19(.A(w2[38]), .B(w2[39]), .Y(w3[19]));
	NAND2_X1A_A12TR level_4_2(.A(w2[4]), .B(w2[5]), .Y(w3[2]));
	NAND2_X1A_A12TR level_4_20(.A(w2[40]), .B(w2[41]), .Y(w3[20]));
	NAND2_X1A_A12TR level_4_21(.A(w2[42]), .B(w2[43]), .Y(w3[21]));
	NAND2_X1A_A12TR level_4_22(.A(w2[44]), .B(w2[45]), .Y(w3[22]));
	NAND2_X1A_A12TR level_4_23(.A(w2[46]), .B(w2[47]), .Y(w3[23]));
	NAND2_X1A_A12TR level_4_24(.A(w2[48]), .B(w2[49]), .Y(w3[24]));
	NAND2_X1A_A12TR level_4_25(.A(w2[50]), .B(w2[51]), .Y(w3[25]));
	NAND2_X1A_A12TR level_4_26(.A(w2[52]), .B(w2[53]), .Y(w3[26]));
	NAND2_X1A_A12TR level_4_27(.A(w2[54]), .B(w2[55]), .Y(w3[27]));
	NAND2_X1A_A12TR level_4_28(.A(w2[56]), .B(w2[57]), .Y(w3[28]));
	NAND2_X1A_A12TR level_4_29(.A(w2[58]), .B(w2[59]), .Y(w3[29]));
	NAND2_X1A_A12TR level_4_3(.A(w2[6]), .B(w2[7]), .Y(w3[3]));
	NAND2_X1A_A12TR level_4_30(.A(w2[60]), .B(w2[61]), .Y(w3[30]));
	NAND2_X1A_A12TR level_4_31(.A(w2[62]), .B(w2[63]), .Y(w3[31]));
	NAND2_X1A_A12TR level_4_4(.A(w2[8]), .B(w2[9]), .Y(w3[4]));
	NAND2_X1A_A12TR level_4_5(.A(w2[10]), .B(w2[11]), .Y(w3[5]));
	NAND2_X1A_A12TR level_4_6(.A(w2[12]), .B(w2[13]), .Y(w3[6]));
	NAND2_X1A_A12TR level_4_7(.A(w2[14]), .B(w2[15]), .Y(w3[7]));
	NAND2_X1A_A12TR level_4_8(.A(w2[16]), .B(w2[17]), .Y(w3[8]));
	NAND2_X1A_A12TR level_4_9(.A(w2[18]), .B(w2[19]), .Y(w3[9]));
	NOR2_X1A_A12TR level_5_0(.A(w3[0]), .B(w3[1]), .Y(w4[0]));
	NOR2_X1A_A12TR level_5_1(.A(w3[2]), .B(w3[3]), .Y(w4[1]));
	NOR2_X1A_A12TR level_5_10(.A(w3[20]), .B(w3[21]), .Y(w4[10]));
	NOR2_X1A_A12TR level_5_11(.A(w3[22]), .B(w3[23]), .Y(w4[11]));
	NOR2_X1A_A12TR level_5_12(.A(w3[24]), .B(w3[25]), .Y(w4[12]));
	NOR2_X1A_A12TR level_5_13(.A(w3[26]), .B(w3[27]), .Y(w4[13]));
	NOR2_X1A_A12TR level_5_14(.A(w3[28]), .B(w3[29]), .Y(w4[14]));
	NOR2_X1A_A12TR level_5_15(.A(w3[30]), .B(w3[31]), .Y(w4[15]));
	NOR2_X1A_A12TR level_5_2(.A(w3[4]), .B(w3[5]), .Y(w4[2]));
	NOR2_X1A_A12TR level_5_3(.A(w3[6]), .B(w3[7]), .Y(w4[3]));
	NOR2_X1A_A12TR level_5_4(.A(w3[8]), .B(w3[9]), .Y(w4[4]));
	NOR2_X1A_A12TR level_5_5(.A(w3[10]), .B(w3[11]), .Y(w4[5]));
	NOR2_X1A_A12TR level_5_6(.A(w3[12]), .B(w3[13]), .Y(w4[6]));
	NOR2_X1A_A12TR level_5_7(.A(w3[14]), .B(w3[15]), .Y(w4[7]));
	NOR2_X1A_A12TR level_5_8(.A(w3[16]), .B(w3[17]), .Y(w4[8]));
	NOR2_X1A_A12TR level_5_9(.A(w3[18]), .B(w3[19]), .Y(w4[9]));
	NAND2_X1A_A12TR level_6_0(.A(w4[0]), .B(w4[1]), .Y(w5[0]));
	NAND2_X1A_A12TR level_6_1(.A(w4[2]), .B(w4[3]), .Y(w5[1]));
	NAND2_X1A_A12TR level_6_2(.A(w4[4]), .B(w4[5]), .Y(w5[2]));
	NAND2_X1A_A12TR level_6_3(.A(w4[6]), .B(w4[7]), .Y(w5[3]));
	NAND2_X1A_A12TR level_6_4(.A(w4[8]), .B(w4[9]), .Y(w5[4]));
	NAND2_X1A_A12TR level_6_5(.A(w4[10]), .B(w4[11]), .Y(w5[5]));
	NAND2_X1A_A12TR level_6_6(.A(w4[12]), .B(w4[13]), .Y(w5[6]));
	NAND2_X1A_A12TR level_6_7(.A(w4[14]), .B(w4[15]), .Y(w5[7]));
	NOR2_X1A_A12TR level_7_0(.A(w5[0]), .B(w5[1]), .Y(w6[0]));
	NOR2_X1A_A12TR level_7_1(.A(w5[2]), .B(w5[3]), .Y(w6[1]));
	NOR2_X1A_A12TR level_7_2(.A(w5[4]), .B(w5[5]), .Y(w6[2]));
	NOR2_X1A_A12TR level_7_3(.A(w5[6]), .B(w5[7]), .Y(w6[3]));
	NAND2_X1A_A12TR level_8_0(.A(w6[0]), .B(w6[1]), .Y(w7[0]));
	NAND2_X1A_A12TR level_8_1(.A(w6[2]), .B(w6[3]), .Y(w7[1]));
	NOR2_X1A_A12TR level_9_0(.A(w7[0]), .B(w7[1]), .Y(w8[0]));

endmodule
