

module rwlBuff_strip (IN, OUT);

	//ports
	output [255:0] OUT;
	input [255:0] IN;

	//wires
	wire [255:0] OUT;
	wire [255:0] IN;

	//instances
	BUFH_X3M_A12TR rwlBuff_0(.A(IN[0]), .Y(OUT[0]));
	BUFH_X3M_A12TR rwlBuff_1(.A(IN[1]), .Y(OUT[1]));
	BUFH_X3M_A12TR rwlBuff_10(.A(IN[10]), .Y(OUT[10]));
	BUFH_X3M_A12TR rwlBuff_100(.A(IN[100]), .Y(OUT[100]));
	BUFH_X3M_A12TR rwlBuff_101(.A(IN[101]), .Y(OUT[101]));
	BUFH_X3M_A12TR rwlBuff_102(.A(IN[102]), .Y(OUT[102]));
	BUFH_X3M_A12TR rwlBuff_103(.A(IN[103]), .Y(OUT[103]));
	BUFH_X3M_A12TR rwlBuff_104(.A(IN[104]), .Y(OUT[104]));
	BUFH_X3M_A12TR rwlBuff_105(.A(IN[105]), .Y(OUT[105]));
	BUFH_X3M_A12TR rwlBuff_106(.A(IN[106]), .Y(OUT[106]));
	BUFH_X3M_A12TR rwlBuff_107(.A(IN[107]), .Y(OUT[107]));
	BUFH_X3M_A12TR rwlBuff_108(.A(IN[108]), .Y(OUT[108]));
	BUFH_X3M_A12TR rwlBuff_109(.A(IN[109]), .Y(OUT[109]));
	BUFH_X3M_A12TR rwlBuff_11(.A(IN[11]), .Y(OUT[11]));
	BUFH_X3M_A12TR rwlBuff_110(.A(IN[110]), .Y(OUT[110]));
	BUFH_X3M_A12TR rwlBuff_111(.A(IN[111]), .Y(OUT[111]));
	BUFH_X3M_A12TR rwlBuff_112(.A(IN[112]), .Y(OUT[112]));
	BUFH_X3M_A12TR rwlBuff_113(.A(IN[113]), .Y(OUT[113]));
	BUFH_X3M_A12TR rwlBuff_114(.A(IN[114]), .Y(OUT[114]));
	BUFH_X3M_A12TR rwlBuff_115(.A(IN[115]), .Y(OUT[115]));
	BUFH_X3M_A12TR rwlBuff_116(.A(IN[116]), .Y(OUT[116]));
	BUFH_X3M_A12TR rwlBuff_117(.A(IN[117]), .Y(OUT[117]));
	BUFH_X3M_A12TR rwlBuff_118(.A(IN[118]), .Y(OUT[118]));
	BUFH_X3M_A12TR rwlBuff_119(.A(IN[119]), .Y(OUT[119]));
	BUFH_X3M_A12TR rwlBuff_12(.A(IN[12]), .Y(OUT[12]));
	BUFH_X3M_A12TR rwlBuff_120(.A(IN[120]), .Y(OUT[120]));
	BUFH_X3M_A12TR rwlBuff_121(.A(IN[121]), .Y(OUT[121]));
	BUFH_X3M_A12TR rwlBuff_122(.A(IN[122]), .Y(OUT[122]));
	BUFH_X3M_A12TR rwlBuff_123(.A(IN[123]), .Y(OUT[123]));
	BUFH_X3M_A12TR rwlBuff_124(.A(IN[124]), .Y(OUT[124]));
	BUFH_X3M_A12TR rwlBuff_125(.A(IN[125]), .Y(OUT[125]));
	BUFH_X3M_A12TR rwlBuff_126(.A(IN[126]), .Y(OUT[126]));
	BUFH_X3M_A12TR rwlBuff_127(.A(IN[127]), .Y(OUT[127]));
	BUFH_X3M_A12TR rwlBuff_128(.A(IN[128]), .Y(OUT[128]));
	BUFH_X3M_A12TR rwlBuff_129(.A(IN[129]), .Y(OUT[129]));
	BUFH_X3M_A12TR rwlBuff_13(.A(IN[13]), .Y(OUT[13]));
	BUFH_X3M_A12TR rwlBuff_130(.A(IN[130]), .Y(OUT[130]));
	BUFH_X3M_A12TR rwlBuff_131(.A(IN[131]), .Y(OUT[131]));
	BUFH_X3M_A12TR rwlBuff_132(.A(IN[132]), .Y(OUT[132]));
	BUFH_X3M_A12TR rwlBuff_133(.A(IN[133]), .Y(OUT[133]));
	BUFH_X3M_A12TR rwlBuff_134(.A(IN[134]), .Y(OUT[134]));
	BUFH_X3M_A12TR rwlBuff_135(.A(IN[135]), .Y(OUT[135]));
	BUFH_X3M_A12TR rwlBuff_136(.A(IN[136]), .Y(OUT[136]));
	BUFH_X3M_A12TR rwlBuff_137(.A(IN[137]), .Y(OUT[137]));
	BUFH_X3M_A12TR rwlBuff_138(.A(IN[138]), .Y(OUT[138]));
	BUFH_X3M_A12TR rwlBuff_139(.A(IN[139]), .Y(OUT[139]));
	BUFH_X3M_A12TR rwlBuff_14(.A(IN[14]), .Y(OUT[14]));
	BUFH_X3M_A12TR rwlBuff_140(.A(IN[140]), .Y(OUT[140]));
	BUFH_X3M_A12TR rwlBuff_141(.A(IN[141]), .Y(OUT[141]));
	BUFH_X3M_A12TR rwlBuff_142(.A(IN[142]), .Y(OUT[142]));
	BUFH_X3M_A12TR rwlBuff_143(.A(IN[143]), .Y(OUT[143]));
	BUFH_X3M_A12TR rwlBuff_144(.A(IN[144]), .Y(OUT[144]));
	BUFH_X3M_A12TR rwlBuff_145(.A(IN[145]), .Y(OUT[145]));
	BUFH_X3M_A12TR rwlBuff_146(.A(IN[146]), .Y(OUT[146]));
	BUFH_X3M_A12TR rwlBuff_147(.A(IN[147]), .Y(OUT[147]));
	BUFH_X3M_A12TR rwlBuff_148(.A(IN[148]), .Y(OUT[148]));
	BUFH_X3M_A12TR rwlBuff_149(.A(IN[149]), .Y(OUT[149]));
	BUFH_X3M_A12TR rwlBuff_15(.A(IN[15]), .Y(OUT[15]));
	BUFH_X3M_A12TR rwlBuff_150(.A(IN[150]), .Y(OUT[150]));
	BUFH_X3M_A12TR rwlBuff_151(.A(IN[151]), .Y(OUT[151]));
	BUFH_X3M_A12TR rwlBuff_152(.A(IN[152]), .Y(OUT[152]));
	BUFH_X3M_A12TR rwlBuff_153(.A(IN[153]), .Y(OUT[153]));
	BUFH_X3M_A12TR rwlBuff_154(.A(IN[154]), .Y(OUT[154]));
	BUFH_X3M_A12TR rwlBuff_155(.A(IN[155]), .Y(OUT[155]));
	BUFH_X3M_A12TR rwlBuff_156(.A(IN[156]), .Y(OUT[156]));
	BUFH_X3M_A12TR rwlBuff_157(.A(IN[157]), .Y(OUT[157]));
	BUFH_X3M_A12TR rwlBuff_158(.A(IN[158]), .Y(OUT[158]));
	BUFH_X3M_A12TR rwlBuff_159(.A(IN[159]), .Y(OUT[159]));
	BUFH_X3M_A12TR rwlBuff_16(.A(IN[16]), .Y(OUT[16]));
	BUFH_X3M_A12TR rwlBuff_160(.A(IN[160]), .Y(OUT[160]));
	BUFH_X3M_A12TR rwlBuff_161(.A(IN[161]), .Y(OUT[161]));
	BUFH_X3M_A12TR rwlBuff_162(.A(IN[162]), .Y(OUT[162]));
	BUFH_X3M_A12TR rwlBuff_163(.A(IN[163]), .Y(OUT[163]));
	BUFH_X3M_A12TR rwlBuff_164(.A(IN[164]), .Y(OUT[164]));
	BUFH_X3M_A12TR rwlBuff_165(.A(IN[165]), .Y(OUT[165]));
	BUFH_X3M_A12TR rwlBuff_166(.A(IN[166]), .Y(OUT[166]));
	BUFH_X3M_A12TR rwlBuff_167(.A(IN[167]), .Y(OUT[167]));
	BUFH_X3M_A12TR rwlBuff_168(.A(IN[168]), .Y(OUT[168]));
	BUFH_X3M_A12TR rwlBuff_169(.A(IN[169]), .Y(OUT[169]));
	BUFH_X3M_A12TR rwlBuff_17(.A(IN[17]), .Y(OUT[17]));
	BUFH_X3M_A12TR rwlBuff_170(.A(IN[170]), .Y(OUT[170]));
	BUFH_X3M_A12TR rwlBuff_171(.A(IN[171]), .Y(OUT[171]));
	BUFH_X3M_A12TR rwlBuff_172(.A(IN[172]), .Y(OUT[172]));
	BUFH_X3M_A12TR rwlBuff_173(.A(IN[173]), .Y(OUT[173]));
	BUFH_X3M_A12TR rwlBuff_174(.A(IN[174]), .Y(OUT[174]));
	BUFH_X3M_A12TR rwlBuff_175(.A(IN[175]), .Y(OUT[175]));
	BUFH_X3M_A12TR rwlBuff_176(.A(IN[176]), .Y(OUT[176]));
	BUFH_X3M_A12TR rwlBuff_177(.A(IN[177]), .Y(OUT[177]));
	BUFH_X3M_A12TR rwlBuff_178(.A(IN[178]), .Y(OUT[178]));
	BUFH_X3M_A12TR rwlBuff_179(.A(IN[179]), .Y(OUT[179]));
	BUFH_X3M_A12TR rwlBuff_18(.A(IN[18]), .Y(OUT[18]));
	BUFH_X3M_A12TR rwlBuff_180(.A(IN[180]), .Y(OUT[180]));
	BUFH_X3M_A12TR rwlBuff_181(.A(IN[181]), .Y(OUT[181]));
	BUFH_X3M_A12TR rwlBuff_182(.A(IN[182]), .Y(OUT[182]));
	BUFH_X3M_A12TR rwlBuff_183(.A(IN[183]), .Y(OUT[183]));
	BUFH_X3M_A12TR rwlBuff_184(.A(IN[184]), .Y(OUT[184]));
	BUFH_X3M_A12TR rwlBuff_185(.A(IN[185]), .Y(OUT[185]));
	BUFH_X3M_A12TR rwlBuff_186(.A(IN[186]), .Y(OUT[186]));
	BUFH_X3M_A12TR rwlBuff_187(.A(IN[187]), .Y(OUT[187]));
	BUFH_X3M_A12TR rwlBuff_188(.A(IN[188]), .Y(OUT[188]));
	BUFH_X3M_A12TR rwlBuff_189(.A(IN[189]), .Y(OUT[189]));
	BUFH_X3M_A12TR rwlBuff_19(.A(IN[19]), .Y(OUT[19]));
	BUFH_X3M_A12TR rwlBuff_190(.A(IN[190]), .Y(OUT[190]));
	BUFH_X3M_A12TR rwlBuff_191(.A(IN[191]), .Y(OUT[191]));
	BUFH_X3M_A12TR rwlBuff_192(.A(IN[192]), .Y(OUT[192]));
	BUFH_X3M_A12TR rwlBuff_193(.A(IN[193]), .Y(OUT[193]));
	BUFH_X3M_A12TR rwlBuff_194(.A(IN[194]), .Y(OUT[194]));
	BUFH_X3M_A12TR rwlBuff_195(.A(IN[195]), .Y(OUT[195]));
	BUFH_X3M_A12TR rwlBuff_196(.A(IN[196]), .Y(OUT[196]));
	BUFH_X3M_A12TR rwlBuff_197(.A(IN[197]), .Y(OUT[197]));
	BUFH_X3M_A12TR rwlBuff_198(.A(IN[198]), .Y(OUT[198]));
	BUFH_X3M_A12TR rwlBuff_199(.A(IN[199]), .Y(OUT[199]));
	BUFH_X3M_A12TR rwlBuff_2(.A(IN[2]), .Y(OUT[2]));
	BUFH_X3M_A12TR rwlBuff_20(.A(IN[20]), .Y(OUT[20]));
	BUFH_X3M_A12TR rwlBuff_200(.A(IN[200]), .Y(OUT[200]));
	BUFH_X3M_A12TR rwlBuff_201(.A(IN[201]), .Y(OUT[201]));
	BUFH_X3M_A12TR rwlBuff_202(.A(IN[202]), .Y(OUT[202]));
	BUFH_X3M_A12TR rwlBuff_203(.A(IN[203]), .Y(OUT[203]));
	BUFH_X3M_A12TR rwlBuff_204(.A(IN[204]), .Y(OUT[204]));
	BUFH_X3M_A12TR rwlBuff_205(.A(IN[205]), .Y(OUT[205]));
	BUFH_X3M_A12TR rwlBuff_206(.A(IN[206]), .Y(OUT[206]));
	BUFH_X3M_A12TR rwlBuff_207(.A(IN[207]), .Y(OUT[207]));
	BUFH_X3M_A12TR rwlBuff_208(.A(IN[208]), .Y(OUT[208]));
	BUFH_X3M_A12TR rwlBuff_209(.A(IN[209]), .Y(OUT[209]));
	BUFH_X3M_A12TR rwlBuff_21(.A(IN[21]), .Y(OUT[21]));
	BUFH_X3M_A12TR rwlBuff_210(.A(IN[210]), .Y(OUT[210]));
	BUFH_X3M_A12TR rwlBuff_211(.A(IN[211]), .Y(OUT[211]));
	BUFH_X3M_A12TR rwlBuff_212(.A(IN[212]), .Y(OUT[212]));
	BUFH_X3M_A12TR rwlBuff_213(.A(IN[213]), .Y(OUT[213]));
	BUFH_X3M_A12TR rwlBuff_214(.A(IN[214]), .Y(OUT[214]));
	BUFH_X3M_A12TR rwlBuff_215(.A(IN[215]), .Y(OUT[215]));
	BUFH_X3M_A12TR rwlBuff_216(.A(IN[216]), .Y(OUT[216]));
	BUFH_X3M_A12TR rwlBuff_217(.A(IN[217]), .Y(OUT[217]));
	BUFH_X3M_A12TR rwlBuff_218(.A(IN[218]), .Y(OUT[218]));
	BUFH_X3M_A12TR rwlBuff_219(.A(IN[219]), .Y(OUT[219]));
	BUFH_X3M_A12TR rwlBuff_22(.A(IN[22]), .Y(OUT[22]));
	BUFH_X3M_A12TR rwlBuff_220(.A(IN[220]), .Y(OUT[220]));
	BUFH_X3M_A12TR rwlBuff_221(.A(IN[221]), .Y(OUT[221]));
	BUFH_X3M_A12TR rwlBuff_222(.A(IN[222]), .Y(OUT[222]));
	BUFH_X3M_A12TR rwlBuff_223(.A(IN[223]), .Y(OUT[223]));
	BUFH_X3M_A12TR rwlBuff_224(.A(IN[224]), .Y(OUT[224]));
	BUFH_X3M_A12TR rwlBuff_225(.A(IN[225]), .Y(OUT[225]));
	BUFH_X3M_A12TR rwlBuff_226(.A(IN[226]), .Y(OUT[226]));
	BUFH_X3M_A12TR rwlBuff_227(.A(IN[227]), .Y(OUT[227]));
	BUFH_X3M_A12TR rwlBuff_228(.A(IN[228]), .Y(OUT[228]));
	BUFH_X3M_A12TR rwlBuff_229(.A(IN[229]), .Y(OUT[229]));
	BUFH_X3M_A12TR rwlBuff_23(.A(IN[23]), .Y(OUT[23]));
	BUFH_X3M_A12TR rwlBuff_230(.A(IN[230]), .Y(OUT[230]));
	BUFH_X3M_A12TR rwlBuff_231(.A(IN[231]), .Y(OUT[231]));
	BUFH_X3M_A12TR rwlBuff_232(.A(IN[232]), .Y(OUT[232]));
	BUFH_X3M_A12TR rwlBuff_233(.A(IN[233]), .Y(OUT[233]));
	BUFH_X3M_A12TR rwlBuff_234(.A(IN[234]), .Y(OUT[234]));
	BUFH_X3M_A12TR rwlBuff_235(.A(IN[235]), .Y(OUT[235]));
	BUFH_X3M_A12TR rwlBuff_236(.A(IN[236]), .Y(OUT[236]));
	BUFH_X3M_A12TR rwlBuff_237(.A(IN[237]), .Y(OUT[237]));
	BUFH_X3M_A12TR rwlBuff_238(.A(IN[238]), .Y(OUT[238]));
	BUFH_X3M_A12TR rwlBuff_239(.A(IN[239]), .Y(OUT[239]));
	BUFH_X3M_A12TR rwlBuff_24(.A(IN[24]), .Y(OUT[24]));
	BUFH_X3M_A12TR rwlBuff_240(.A(IN[240]), .Y(OUT[240]));
	BUFH_X3M_A12TR rwlBuff_241(.A(IN[241]), .Y(OUT[241]));
	BUFH_X3M_A12TR rwlBuff_242(.A(IN[242]), .Y(OUT[242]));
	BUFH_X3M_A12TR rwlBuff_243(.A(IN[243]), .Y(OUT[243]));
	BUFH_X3M_A12TR rwlBuff_244(.A(IN[244]), .Y(OUT[244]));
	BUFH_X3M_A12TR rwlBuff_245(.A(IN[245]), .Y(OUT[245]));
	BUFH_X3M_A12TR rwlBuff_246(.A(IN[246]), .Y(OUT[246]));
	BUFH_X3M_A12TR rwlBuff_247(.A(IN[247]), .Y(OUT[247]));
	BUFH_X3M_A12TR rwlBuff_248(.A(IN[248]), .Y(OUT[248]));
	BUFH_X3M_A12TR rwlBuff_249(.A(IN[249]), .Y(OUT[249]));
	BUFH_X3M_A12TR rwlBuff_25(.A(IN[25]), .Y(OUT[25]));
	BUFH_X3M_A12TR rwlBuff_250(.A(IN[250]), .Y(OUT[250]));
	BUFH_X3M_A12TR rwlBuff_251(.A(IN[251]), .Y(OUT[251]));
	BUFH_X3M_A12TR rwlBuff_252(.A(IN[252]), .Y(OUT[252]));
	BUFH_X3M_A12TR rwlBuff_253(.A(IN[253]), .Y(OUT[253]));
	BUFH_X3M_A12TR rwlBuff_254(.A(IN[254]), .Y(OUT[254]));
	BUFH_X3M_A12TR rwlBuff_255(.A(IN[255]), .Y(OUT[255]));
	BUFH_X3M_A12TR rwlBuff_26(.A(IN[26]), .Y(OUT[26]));
	BUFH_X3M_A12TR rwlBuff_27(.A(IN[27]), .Y(OUT[27]));
	BUFH_X3M_A12TR rwlBuff_28(.A(IN[28]), .Y(OUT[28]));
	BUFH_X3M_A12TR rwlBuff_29(.A(IN[29]), .Y(OUT[29]));
	BUFH_X3M_A12TR rwlBuff_3(.A(IN[3]), .Y(OUT[3]));
	BUFH_X3M_A12TR rwlBuff_30(.A(IN[30]), .Y(OUT[30]));
	BUFH_X3M_A12TR rwlBuff_31(.A(IN[31]), .Y(OUT[31]));
	BUFH_X3M_A12TR rwlBuff_32(.A(IN[32]), .Y(OUT[32]));
	BUFH_X3M_A12TR rwlBuff_33(.A(IN[33]), .Y(OUT[33]));
	BUFH_X3M_A12TR rwlBuff_34(.A(IN[34]), .Y(OUT[34]));
	BUFH_X3M_A12TR rwlBuff_35(.A(IN[35]), .Y(OUT[35]));
	BUFH_X3M_A12TR rwlBuff_36(.A(IN[36]), .Y(OUT[36]));
	BUFH_X3M_A12TR rwlBuff_37(.A(IN[37]), .Y(OUT[37]));
	BUFH_X3M_A12TR rwlBuff_38(.A(IN[38]), .Y(OUT[38]));
	BUFH_X3M_A12TR rwlBuff_39(.A(IN[39]), .Y(OUT[39]));
	BUFH_X3M_A12TR rwlBuff_4(.A(IN[4]), .Y(OUT[4]));
	BUFH_X3M_A12TR rwlBuff_40(.A(IN[40]), .Y(OUT[40]));
	BUFH_X3M_A12TR rwlBuff_41(.A(IN[41]), .Y(OUT[41]));
	BUFH_X3M_A12TR rwlBuff_42(.A(IN[42]), .Y(OUT[42]));
	BUFH_X3M_A12TR rwlBuff_43(.A(IN[43]), .Y(OUT[43]));
	BUFH_X3M_A12TR rwlBuff_44(.A(IN[44]), .Y(OUT[44]));
	BUFH_X3M_A12TR rwlBuff_45(.A(IN[45]), .Y(OUT[45]));
	BUFH_X3M_A12TR rwlBuff_46(.A(IN[46]), .Y(OUT[46]));
	BUFH_X3M_A12TR rwlBuff_47(.A(IN[47]), .Y(OUT[47]));
	BUFH_X3M_A12TR rwlBuff_48(.A(IN[48]), .Y(OUT[48]));
	BUFH_X3M_A12TR rwlBuff_49(.A(IN[49]), .Y(OUT[49]));
	BUFH_X3M_A12TR rwlBuff_5(.A(IN[5]), .Y(OUT[5]));
	BUFH_X3M_A12TR rwlBuff_50(.A(IN[50]), .Y(OUT[50]));
	BUFH_X3M_A12TR rwlBuff_51(.A(IN[51]), .Y(OUT[51]));
	BUFH_X3M_A12TR rwlBuff_52(.A(IN[52]), .Y(OUT[52]));
	BUFH_X3M_A12TR rwlBuff_53(.A(IN[53]), .Y(OUT[53]));
	BUFH_X3M_A12TR rwlBuff_54(.A(IN[54]), .Y(OUT[54]));
	BUFH_X3M_A12TR rwlBuff_55(.A(IN[55]), .Y(OUT[55]));
	BUFH_X3M_A12TR rwlBuff_56(.A(IN[56]), .Y(OUT[56]));
	BUFH_X3M_A12TR rwlBuff_57(.A(IN[57]), .Y(OUT[57]));
	BUFH_X3M_A12TR rwlBuff_58(.A(IN[58]), .Y(OUT[58]));
	BUFH_X3M_A12TR rwlBuff_59(.A(IN[59]), .Y(OUT[59]));
	BUFH_X3M_A12TR rwlBuff_6(.A(IN[6]), .Y(OUT[6]));
	BUFH_X3M_A12TR rwlBuff_60(.A(IN[60]), .Y(OUT[60]));
	BUFH_X3M_A12TR rwlBuff_61(.A(IN[61]), .Y(OUT[61]));
	BUFH_X3M_A12TR rwlBuff_62(.A(IN[62]), .Y(OUT[62]));
	BUFH_X3M_A12TR rwlBuff_63(.A(IN[63]), .Y(OUT[63]));
	BUFH_X3M_A12TR rwlBuff_64(.A(IN[64]), .Y(OUT[64]));
	BUFH_X3M_A12TR rwlBuff_65(.A(IN[65]), .Y(OUT[65]));
	BUFH_X3M_A12TR rwlBuff_66(.A(IN[66]), .Y(OUT[66]));
	BUFH_X3M_A12TR rwlBuff_67(.A(IN[67]), .Y(OUT[67]));
	BUFH_X3M_A12TR rwlBuff_68(.A(IN[68]), .Y(OUT[68]));
	BUFH_X3M_A12TR rwlBuff_69(.A(IN[69]), .Y(OUT[69]));
	BUFH_X3M_A12TR rwlBuff_7(.A(IN[7]), .Y(OUT[7]));
	BUFH_X3M_A12TR rwlBuff_70(.A(IN[70]), .Y(OUT[70]));
	BUFH_X3M_A12TR rwlBuff_71(.A(IN[71]), .Y(OUT[71]));
	BUFH_X3M_A12TR rwlBuff_72(.A(IN[72]), .Y(OUT[72]));
	BUFH_X3M_A12TR rwlBuff_73(.A(IN[73]), .Y(OUT[73]));
	BUFH_X3M_A12TR rwlBuff_74(.A(IN[74]), .Y(OUT[74]));
	BUFH_X3M_A12TR rwlBuff_75(.A(IN[75]), .Y(OUT[75]));
	BUFH_X3M_A12TR rwlBuff_76(.A(IN[76]), .Y(OUT[76]));
	BUFH_X3M_A12TR rwlBuff_77(.A(IN[77]), .Y(OUT[77]));
	BUFH_X3M_A12TR rwlBuff_78(.A(IN[78]), .Y(OUT[78]));
	BUFH_X3M_A12TR rwlBuff_79(.A(IN[79]), .Y(OUT[79]));
	BUFH_X3M_A12TR rwlBuff_8(.A(IN[8]), .Y(OUT[8]));
	BUFH_X3M_A12TR rwlBuff_80(.A(IN[80]), .Y(OUT[80]));
	BUFH_X3M_A12TR rwlBuff_81(.A(IN[81]), .Y(OUT[81]));
	BUFH_X3M_A12TR rwlBuff_82(.A(IN[82]), .Y(OUT[82]));
	BUFH_X3M_A12TR rwlBuff_83(.A(IN[83]), .Y(OUT[83]));
	BUFH_X3M_A12TR rwlBuff_84(.A(IN[84]), .Y(OUT[84]));
	BUFH_X3M_A12TR rwlBuff_85(.A(IN[85]), .Y(OUT[85]));
	BUFH_X3M_A12TR rwlBuff_86(.A(IN[86]), .Y(OUT[86]));
	BUFH_X3M_A12TR rwlBuff_87(.A(IN[87]), .Y(OUT[87]));
	BUFH_X3M_A12TR rwlBuff_88(.A(IN[88]), .Y(OUT[88]));
	BUFH_X3M_A12TR rwlBuff_89(.A(IN[89]), .Y(OUT[89]));
	BUFH_X3M_A12TR rwlBuff_9(.A(IN[9]), .Y(OUT[9]));
	BUFH_X3M_A12TR rwlBuff_90(.A(IN[90]), .Y(OUT[90]));
	BUFH_X3M_A12TR rwlBuff_91(.A(IN[91]), .Y(OUT[91]));
	BUFH_X3M_A12TR rwlBuff_92(.A(IN[92]), .Y(OUT[92]));
	BUFH_X3M_A12TR rwlBuff_93(.A(IN[93]), .Y(OUT[93]));
	BUFH_X3M_A12TR rwlBuff_94(.A(IN[94]), .Y(OUT[94]));
	BUFH_X3M_A12TR rwlBuff_95(.A(IN[95]), .Y(OUT[95]));
	BUFH_X3M_A12TR rwlBuff_96(.A(IN[96]), .Y(OUT[96]));
	BUFH_X3M_A12TR rwlBuff_97(.A(IN[97]), .Y(OUT[97]));
	BUFH_X3M_A12TR rwlBuff_98(.A(IN[98]), .Y(OUT[98]));
	BUFH_X3M_A12TR rwlBuff_99(.A(IN[99]), .Y(OUT[99]));

endmodule
