

module Decoder_3_8 (decoder_in, decoder_out);

    //ports
    input [2:0] decoder_in;
    output [7:0] decoder_out;

    //wires
    wire [2:0] decoder_in;
    wire [7:0] decoder_out;

    //instances

endmodule
