

module welltap_strip ();

	//instances
	WELLANTENNATIEPW2_A12TR welltap_0();
	WELLANTENNATIEPW2_A12TR welltap_1();
	WELLANTENNATIEPW2_A12TR welltap_10();
	WELLANTENNATIEPW2_A12TR welltap_100();
	WELLANTENNATIEPW2_A12TR welltap_101();
	WELLANTENNATIEPW2_A12TR welltap_102();
	WELLANTENNATIEPW2_A12TR welltap_103();
	WELLANTENNATIEPW2_A12TR welltap_104();
	WELLANTENNATIEPW2_A12TR welltap_105();
	WELLANTENNATIEPW2_A12TR welltap_106();
	WELLANTENNATIEPW2_A12TR welltap_107();
	WELLANTENNATIEPW2_A12TR welltap_108();
	WELLANTENNATIEPW2_A12TR welltap_109();
	WELLANTENNATIEPW2_A12TR welltap_11();
	WELLANTENNATIEPW2_A12TR welltap_110();
	WELLANTENNATIEPW2_A12TR welltap_111();
	WELLANTENNATIEPW2_A12TR welltap_112();
	WELLANTENNATIEPW2_A12TR welltap_113();
	WELLANTENNATIEPW2_A12TR welltap_114();
	WELLANTENNATIEPW2_A12TR welltap_115();
	WELLANTENNATIEPW2_A12TR welltap_116();
	WELLANTENNATIEPW2_A12TR welltap_117();
	WELLANTENNATIEPW2_A12TR welltap_118();
	WELLANTENNATIEPW2_A12TR welltap_119();
	WELLANTENNATIEPW2_A12TR welltap_12();
	WELLANTENNATIEPW2_A12TR welltap_120();
	WELLANTENNATIEPW2_A12TR welltap_121();
	WELLANTENNATIEPW2_A12TR welltap_122();
	WELLANTENNATIEPW2_A12TR welltap_123();
	WELLANTENNATIEPW2_A12TR welltap_124();
	WELLANTENNATIEPW2_A12TR welltap_125();
	WELLANTENNATIEPW2_A12TR welltap_126();
	WELLANTENNATIEPW2_A12TR welltap_127();
	WELLANTENNATIEPW2_A12TR welltap_128();
	WELLANTENNATIEPW2_A12TR welltap_129();
	WELLANTENNATIEPW2_A12TR welltap_13();
	WELLANTENNATIEPW2_A12TR welltap_130();
	WELLANTENNATIEPW2_A12TR welltap_131();
	WELLANTENNATIEPW2_A12TR welltap_132();
	WELLANTENNATIEPW2_A12TR welltap_133();
	WELLANTENNATIEPW2_A12TR welltap_134();
	WELLANTENNATIEPW2_A12TR welltap_135();
	WELLANTENNATIEPW2_A12TR welltap_136();
	WELLANTENNATIEPW2_A12TR welltap_137();
	WELLANTENNATIEPW2_A12TR welltap_138();
	WELLANTENNATIEPW2_A12TR welltap_139();
	WELLANTENNATIEPW2_A12TR welltap_14();
	WELLANTENNATIEPW2_A12TR welltap_140();
	WELLANTENNATIEPW2_A12TR welltap_141();
	WELLANTENNATIEPW2_A12TR welltap_142();
	WELLANTENNATIEPW2_A12TR welltap_143();
	WELLANTENNATIEPW2_A12TR welltap_144();
	WELLANTENNATIEPW2_A12TR welltap_145();
	WELLANTENNATIEPW2_A12TR welltap_146();
	WELLANTENNATIEPW2_A12TR welltap_147();
	WELLANTENNATIEPW2_A12TR welltap_148();
	WELLANTENNATIEPW2_A12TR welltap_149();
	WELLANTENNATIEPW2_A12TR welltap_15();
	WELLANTENNATIEPW2_A12TR welltap_150();
	WELLANTENNATIEPW2_A12TR welltap_151();
	WELLANTENNATIEPW2_A12TR welltap_152();
	WELLANTENNATIEPW2_A12TR welltap_153();
	WELLANTENNATIEPW2_A12TR welltap_154();
	WELLANTENNATIEPW2_A12TR welltap_155();
	WELLANTENNATIEPW2_A12TR welltap_156();
	WELLANTENNATIEPW2_A12TR welltap_157();
	WELLANTENNATIEPW2_A12TR welltap_158();
	WELLANTENNATIEPW2_A12TR welltap_159();
	WELLANTENNATIEPW2_A12TR welltap_16();
	WELLANTENNATIEPW2_A12TR welltap_160();
	WELLANTENNATIEPW2_A12TR welltap_161();
	WELLANTENNATIEPW2_A12TR welltap_162();
	WELLANTENNATIEPW2_A12TR welltap_163();
	WELLANTENNATIEPW2_A12TR welltap_164();
	WELLANTENNATIEPW2_A12TR welltap_165();
	WELLANTENNATIEPW2_A12TR welltap_166();
	WELLANTENNATIEPW2_A12TR welltap_167();
	WELLANTENNATIEPW2_A12TR welltap_168();
	WELLANTENNATIEPW2_A12TR welltap_169();
	WELLANTENNATIEPW2_A12TR welltap_17();
	WELLANTENNATIEPW2_A12TR welltap_170();
	WELLANTENNATIEPW2_A12TR welltap_171();
	WELLANTENNATIEPW2_A12TR welltap_172();
	WELLANTENNATIEPW2_A12TR welltap_173();
	WELLANTENNATIEPW2_A12TR welltap_174();
	WELLANTENNATIEPW2_A12TR welltap_175();
	WELLANTENNATIEPW2_A12TR welltap_176();
	WELLANTENNATIEPW2_A12TR welltap_177();
	WELLANTENNATIEPW2_A12TR welltap_178();
	WELLANTENNATIEPW2_A12TR welltap_179();
	WELLANTENNATIEPW2_A12TR welltap_18();
	WELLANTENNATIEPW2_A12TR welltap_180();
	WELLANTENNATIEPW2_A12TR welltap_181();
	WELLANTENNATIEPW2_A12TR welltap_182();
	WELLANTENNATIEPW2_A12TR welltap_183();
	WELLANTENNATIEPW2_A12TR welltap_184();
	WELLANTENNATIEPW2_A12TR welltap_185();
	WELLANTENNATIEPW2_A12TR welltap_186();
	WELLANTENNATIEPW2_A12TR welltap_187();
	WELLANTENNATIEPW2_A12TR welltap_188();
	WELLANTENNATIEPW2_A12TR welltap_189();
	WELLANTENNATIEPW2_A12TR welltap_19();
	WELLANTENNATIEPW2_A12TR welltap_190();
	WELLANTENNATIEPW2_A12TR welltap_191();
	WELLANTENNATIEPW2_A12TR welltap_192();
	WELLANTENNATIEPW2_A12TR welltap_193();
	WELLANTENNATIEPW2_A12TR welltap_194();
	WELLANTENNATIEPW2_A12TR welltap_195();
	WELLANTENNATIEPW2_A12TR welltap_196();
	WELLANTENNATIEPW2_A12TR welltap_197();
	WELLANTENNATIEPW2_A12TR welltap_198();
	WELLANTENNATIEPW2_A12TR welltap_199();
	WELLANTENNATIEPW2_A12TR welltap_2();
	WELLANTENNATIEPW2_A12TR welltap_20();
	WELLANTENNATIEPW2_A12TR welltap_200();
	WELLANTENNATIEPW2_A12TR welltap_201();
	WELLANTENNATIEPW2_A12TR welltap_202();
	WELLANTENNATIEPW2_A12TR welltap_203();
	WELLANTENNATIEPW2_A12TR welltap_204();
	WELLANTENNATIEPW2_A12TR welltap_205();
	WELLANTENNATIEPW2_A12TR welltap_206();
	WELLANTENNATIEPW2_A12TR welltap_207();
	WELLANTENNATIEPW2_A12TR welltap_208();
	WELLANTENNATIEPW2_A12TR welltap_209();
	WELLANTENNATIEPW2_A12TR welltap_21();
	WELLANTENNATIEPW2_A12TR welltap_210();
	WELLANTENNATIEPW2_A12TR welltap_211();
	WELLANTENNATIEPW2_A12TR welltap_212();
	WELLANTENNATIEPW2_A12TR welltap_213();
	WELLANTENNATIEPW2_A12TR welltap_214();
	WELLANTENNATIEPW2_A12TR welltap_215();
	WELLANTENNATIEPW2_A12TR welltap_216();
	WELLANTENNATIEPW2_A12TR welltap_217();
	WELLANTENNATIEPW2_A12TR welltap_218();
	WELLANTENNATIEPW2_A12TR welltap_219();
	WELLANTENNATIEPW2_A12TR welltap_22();
	WELLANTENNATIEPW2_A12TR welltap_220();
	WELLANTENNATIEPW2_A12TR welltap_221();
	WELLANTENNATIEPW2_A12TR welltap_222();
	WELLANTENNATIEPW2_A12TR welltap_223();
	WELLANTENNATIEPW2_A12TR welltap_224();
	WELLANTENNATIEPW2_A12TR welltap_225();
	WELLANTENNATIEPW2_A12TR welltap_226();
	WELLANTENNATIEPW2_A12TR welltap_227();
	WELLANTENNATIEPW2_A12TR welltap_228();
	WELLANTENNATIEPW2_A12TR welltap_229();
	WELLANTENNATIEPW2_A12TR welltap_23();
	WELLANTENNATIEPW2_A12TR welltap_230();
	WELLANTENNATIEPW2_A12TR welltap_231();
	WELLANTENNATIEPW2_A12TR welltap_232();
	WELLANTENNATIEPW2_A12TR welltap_233();
	WELLANTENNATIEPW2_A12TR welltap_234();
	WELLANTENNATIEPW2_A12TR welltap_235();
	WELLANTENNATIEPW2_A12TR welltap_236();
	WELLANTENNATIEPW2_A12TR welltap_237();
	WELLANTENNATIEPW2_A12TR welltap_238();
	WELLANTENNATIEPW2_A12TR welltap_239();
	WELLANTENNATIEPW2_A12TR welltap_24();
	WELLANTENNATIEPW2_A12TR welltap_240();
	WELLANTENNATIEPW2_A12TR welltap_241();
	WELLANTENNATIEPW2_A12TR welltap_242();
	WELLANTENNATIEPW2_A12TR welltap_243();
	WELLANTENNATIEPW2_A12TR welltap_244();
	WELLANTENNATIEPW2_A12TR welltap_245();
	WELLANTENNATIEPW2_A12TR welltap_246();
	WELLANTENNATIEPW2_A12TR welltap_247();
	WELLANTENNATIEPW2_A12TR welltap_248();
	WELLANTENNATIEPW2_A12TR welltap_249();
	WELLANTENNATIEPW2_A12TR welltap_25();
	WELLANTENNATIEPW2_A12TR welltap_250();
	WELLANTENNATIEPW2_A12TR welltap_251();
	WELLANTENNATIEPW2_A12TR welltap_252();
	WELLANTENNATIEPW2_A12TR welltap_253();
	WELLANTENNATIEPW2_A12TR welltap_254();
	WELLANTENNATIEPW2_A12TR welltap_255();
	WELLANTENNATIEPW2_A12TR welltap_256();
	WELLANTENNATIEPW2_A12TR welltap_257();
	WELLANTENNATIEPW2_A12TR welltap_26();
	WELLANTENNATIEPW2_A12TR welltap_27();
	WELLANTENNATIEPW2_A12TR welltap_28();
	WELLANTENNATIEPW2_A12TR welltap_29();
	WELLANTENNATIEPW2_A12TR welltap_3();
	WELLANTENNATIEPW2_A12TR welltap_30();
	WELLANTENNATIEPW2_A12TR welltap_31();
	WELLANTENNATIEPW2_A12TR welltap_32();
	WELLANTENNATIEPW2_A12TR welltap_33();
	WELLANTENNATIEPW2_A12TR welltap_34();
	WELLANTENNATIEPW2_A12TR welltap_35();
	WELLANTENNATIEPW2_A12TR welltap_36();
	WELLANTENNATIEPW2_A12TR welltap_37();
	WELLANTENNATIEPW2_A12TR welltap_38();
	WELLANTENNATIEPW2_A12TR welltap_39();
	WELLANTENNATIEPW2_A12TR welltap_4();
	WELLANTENNATIEPW2_A12TR welltap_40();
	WELLANTENNATIEPW2_A12TR welltap_41();
	WELLANTENNATIEPW2_A12TR welltap_42();
	WELLANTENNATIEPW2_A12TR welltap_43();
	WELLANTENNATIEPW2_A12TR welltap_44();
	WELLANTENNATIEPW2_A12TR welltap_45();
	WELLANTENNATIEPW2_A12TR welltap_46();
	WELLANTENNATIEPW2_A12TR welltap_47();
	WELLANTENNATIEPW2_A12TR welltap_48();
	WELLANTENNATIEPW2_A12TR welltap_49();
	WELLANTENNATIEPW2_A12TR welltap_5();
	WELLANTENNATIEPW2_A12TR welltap_50();
	WELLANTENNATIEPW2_A12TR welltap_51();
	WELLANTENNATIEPW2_A12TR welltap_52();
	WELLANTENNATIEPW2_A12TR welltap_53();
	WELLANTENNATIEPW2_A12TR welltap_54();
	WELLANTENNATIEPW2_A12TR welltap_55();
	WELLANTENNATIEPW2_A12TR welltap_56();
	WELLANTENNATIEPW2_A12TR welltap_57();
	WELLANTENNATIEPW2_A12TR welltap_58();
	WELLANTENNATIEPW2_A12TR welltap_59();
	WELLANTENNATIEPW2_A12TR welltap_6();
	WELLANTENNATIEPW2_A12TR welltap_60();
	WELLANTENNATIEPW2_A12TR welltap_61();
	WELLANTENNATIEPW2_A12TR welltap_62();
	WELLANTENNATIEPW2_A12TR welltap_63();
	WELLANTENNATIEPW2_A12TR welltap_64();
	WELLANTENNATIEPW2_A12TR welltap_65();
	WELLANTENNATIEPW2_A12TR welltap_66();
	WELLANTENNATIEPW2_A12TR welltap_67();
	WELLANTENNATIEPW2_A12TR welltap_68();
	WELLANTENNATIEPW2_A12TR welltap_69();
	WELLANTENNATIEPW2_A12TR welltap_7();
	WELLANTENNATIEPW2_A12TR welltap_70();
	WELLANTENNATIEPW2_A12TR welltap_71();
	WELLANTENNATIEPW2_A12TR welltap_72();
	WELLANTENNATIEPW2_A12TR welltap_73();
	WELLANTENNATIEPW2_A12TR welltap_74();
	WELLANTENNATIEPW2_A12TR welltap_75();
	WELLANTENNATIEPW2_A12TR welltap_76();
	WELLANTENNATIEPW2_A12TR welltap_77();
	WELLANTENNATIEPW2_A12TR welltap_78();
	WELLANTENNATIEPW2_A12TR welltap_79();
	WELLANTENNATIEPW2_A12TR welltap_8();
	WELLANTENNATIEPW2_A12TR welltap_80();
	WELLANTENNATIEPW2_A12TR welltap_81();
	WELLANTENNATIEPW2_A12TR welltap_82();
	WELLANTENNATIEPW2_A12TR welltap_83();
	WELLANTENNATIEPW2_A12TR welltap_84();
	WELLANTENNATIEPW2_A12TR welltap_85();
	WELLANTENNATIEPW2_A12TR welltap_86();
	WELLANTENNATIEPW2_A12TR welltap_87();
	WELLANTENNATIEPW2_A12TR welltap_88();
	WELLANTENNATIEPW2_A12TR welltap_89();
	WELLANTENNATIEPW2_A12TR welltap_9();
	WELLANTENNATIEPW2_A12TR welltap_90();
	WELLANTENNATIEPW2_A12TR welltap_91();
	WELLANTENNATIEPW2_A12TR welltap_92();
	WELLANTENNATIEPW2_A12TR welltap_93();
	WELLANTENNATIEPW2_A12TR welltap_94();
	WELLANTENNATIEPW2_A12TR welltap_95();
	WELLANTENNATIEPW2_A12TR welltap_96();
	WELLANTENNATIEPW2_A12TR welltap_97();
	WELLANTENNATIEPW2_A12TR welltap_98();
	WELLANTENNATIEPW2_A12TR welltap_99();

endmodule
