

module bitslice (DGWCLK, DIN, DOUT, RWL, clk);

	//ports
	input [255:0] RWL;
	input DIN;
	input clk;
	output DOUT;
	input [255:0] DGWCLK;

	//wires
	wire [255:0] RWL;
	wire GDIN;
	wire [255:0] MemoryLatch;
	wire DIN;
	wire clk;
	wire DOUT;
	wire [255:0] DGWCLK;

	//instances
	DFFQ_X2M_A12TR GDIN_reg(.CK(clk), .D(DIN), .Q(GDIN));
	LATQ_X1M_A12TR MemoryLatch_reg_0(.D(GDIN), .G(DGWCLK[0]), .Q(MemoryLatch[0]));
	LATQ_X1M_A12TR MemoryLatch_reg_1(.D(GDIN), .G(DGWCLK[1]), .Q(MemoryLatch[1]));
	LATQ_X1M_A12TR MemoryLatch_reg_10(.D(GDIN), .G(DGWCLK[10]), .Q(MemoryLatch[10]));
	LATQ_X1M_A12TR MemoryLatch_reg_100(.D(GDIN), .G(DGWCLK[100]), .Q(MemoryLatch[100]));
	LATQ_X1M_A12TR MemoryLatch_reg_101(.D(GDIN), .G(DGWCLK[101]), .Q(MemoryLatch[101]));
	LATQ_X1M_A12TR MemoryLatch_reg_102(.D(GDIN), .G(DGWCLK[102]), .Q(MemoryLatch[102]));
	LATQ_X1M_A12TR MemoryLatch_reg_103(.D(GDIN), .G(DGWCLK[103]), .Q(MemoryLatch[103]));
	LATQ_X1M_A12TR MemoryLatch_reg_104(.D(GDIN), .G(DGWCLK[104]), .Q(MemoryLatch[104]));
	LATQ_X1M_A12TR MemoryLatch_reg_105(.D(GDIN), .G(DGWCLK[105]), .Q(MemoryLatch[105]));
	LATQ_X1M_A12TR MemoryLatch_reg_106(.D(GDIN), .G(DGWCLK[106]), .Q(MemoryLatch[106]));
	LATQ_X1M_A12TR MemoryLatch_reg_107(.D(GDIN), .G(DGWCLK[107]), .Q(MemoryLatch[107]));
	LATQ_X1M_A12TR MemoryLatch_reg_108(.D(GDIN), .G(DGWCLK[108]), .Q(MemoryLatch[108]));
	LATQ_X1M_A12TR MemoryLatch_reg_109(.D(GDIN), .G(DGWCLK[109]), .Q(MemoryLatch[109]));
	LATQ_X1M_A12TR MemoryLatch_reg_11(.D(GDIN), .G(DGWCLK[11]), .Q(MemoryLatch[11]));
	LATQ_X1M_A12TR MemoryLatch_reg_110(.D(GDIN), .G(DGWCLK[110]), .Q(MemoryLatch[110]));
	LATQ_X1M_A12TR MemoryLatch_reg_111(.D(GDIN), .G(DGWCLK[111]), .Q(MemoryLatch[111]));
	LATQ_X1M_A12TR MemoryLatch_reg_112(.D(GDIN), .G(DGWCLK[112]), .Q(MemoryLatch[112]));
	LATQ_X1M_A12TR MemoryLatch_reg_113(.D(GDIN), .G(DGWCLK[113]), .Q(MemoryLatch[113]));
	LATQ_X1M_A12TR MemoryLatch_reg_114(.D(GDIN), .G(DGWCLK[114]), .Q(MemoryLatch[114]));
	LATQ_X1M_A12TR MemoryLatch_reg_115(.D(GDIN), .G(DGWCLK[115]), .Q(MemoryLatch[115]));
	LATQ_X1M_A12TR MemoryLatch_reg_116(.D(GDIN), .G(DGWCLK[116]), .Q(MemoryLatch[116]));
	LATQ_X1M_A12TR MemoryLatch_reg_117(.D(GDIN), .G(DGWCLK[117]), .Q(MemoryLatch[117]));
	LATQ_X1M_A12TR MemoryLatch_reg_118(.D(GDIN), .G(DGWCLK[118]), .Q(MemoryLatch[118]));
	LATQ_X1M_A12TR MemoryLatch_reg_119(.D(GDIN), .G(DGWCLK[119]), .Q(MemoryLatch[119]));
	LATQ_X1M_A12TR MemoryLatch_reg_12(.D(GDIN), .G(DGWCLK[12]), .Q(MemoryLatch[12]));
	LATQ_X1M_A12TR MemoryLatch_reg_120(.D(GDIN), .G(DGWCLK[120]), .Q(MemoryLatch[120]));
	LATQ_X1M_A12TR MemoryLatch_reg_121(.D(GDIN), .G(DGWCLK[121]), .Q(MemoryLatch[121]));
	LATQ_X1M_A12TR MemoryLatch_reg_122(.D(GDIN), .G(DGWCLK[122]), .Q(MemoryLatch[122]));
	LATQ_X1M_A12TR MemoryLatch_reg_123(.D(GDIN), .G(DGWCLK[123]), .Q(MemoryLatch[123]));
	LATQ_X1M_A12TR MemoryLatch_reg_124(.D(GDIN), .G(DGWCLK[124]), .Q(MemoryLatch[124]));
	LATQ_X1M_A12TR MemoryLatch_reg_125(.D(GDIN), .G(DGWCLK[125]), .Q(MemoryLatch[125]));
	LATQ_X1M_A12TR MemoryLatch_reg_126(.D(GDIN), .G(DGWCLK[126]), .Q(MemoryLatch[126]));
	LATQ_X1M_A12TR MemoryLatch_reg_127(.D(GDIN), .G(DGWCLK[127]), .Q(MemoryLatch[127]));
	LATQ_X1M_A12TR MemoryLatch_reg_128(.D(GDIN), .G(DGWCLK[128]), .Q(MemoryLatch[128]));
	LATQ_X1M_A12TR MemoryLatch_reg_129(.D(GDIN), .G(DGWCLK[129]), .Q(MemoryLatch[129]));
	LATQ_X1M_A12TR MemoryLatch_reg_13(.D(GDIN), .G(DGWCLK[13]), .Q(MemoryLatch[13]));
	LATQ_X1M_A12TR MemoryLatch_reg_130(.D(GDIN), .G(DGWCLK[130]), .Q(MemoryLatch[130]));
	LATQ_X1M_A12TR MemoryLatch_reg_131(.D(GDIN), .G(DGWCLK[131]), .Q(MemoryLatch[131]));
	LATQ_X1M_A12TR MemoryLatch_reg_132(.D(GDIN), .G(DGWCLK[132]), .Q(MemoryLatch[132]));
	LATQ_X1M_A12TR MemoryLatch_reg_133(.D(GDIN), .G(DGWCLK[133]), .Q(MemoryLatch[133]));
	LATQ_X1M_A12TR MemoryLatch_reg_134(.D(GDIN), .G(DGWCLK[134]), .Q(MemoryLatch[134]));
	LATQ_X1M_A12TR MemoryLatch_reg_135(.D(GDIN), .G(DGWCLK[135]), .Q(MemoryLatch[135]));
	LATQ_X1M_A12TR MemoryLatch_reg_136(.D(GDIN), .G(DGWCLK[136]), .Q(MemoryLatch[136]));
	LATQ_X1M_A12TR MemoryLatch_reg_137(.D(GDIN), .G(DGWCLK[137]), .Q(MemoryLatch[137]));
	LATQ_X1M_A12TR MemoryLatch_reg_138(.D(GDIN), .G(DGWCLK[138]), .Q(MemoryLatch[138]));
	LATQ_X1M_A12TR MemoryLatch_reg_139(.D(GDIN), .G(DGWCLK[139]), .Q(MemoryLatch[139]));
	LATQ_X1M_A12TR MemoryLatch_reg_14(.D(GDIN), .G(DGWCLK[14]), .Q(MemoryLatch[14]));
	LATQ_X1M_A12TR MemoryLatch_reg_140(.D(GDIN), .G(DGWCLK[140]), .Q(MemoryLatch[140]));
	LATQ_X1M_A12TR MemoryLatch_reg_141(.D(GDIN), .G(DGWCLK[141]), .Q(MemoryLatch[141]));
	LATQ_X1M_A12TR MemoryLatch_reg_142(.D(GDIN), .G(DGWCLK[142]), .Q(MemoryLatch[142]));
	LATQ_X1M_A12TR MemoryLatch_reg_143(.D(GDIN), .G(DGWCLK[143]), .Q(MemoryLatch[143]));
	LATQ_X1M_A12TR MemoryLatch_reg_144(.D(GDIN), .G(DGWCLK[144]), .Q(MemoryLatch[144]));
	LATQ_X1M_A12TR MemoryLatch_reg_145(.D(GDIN), .G(DGWCLK[145]), .Q(MemoryLatch[145]));
	LATQ_X1M_A12TR MemoryLatch_reg_146(.D(GDIN), .G(DGWCLK[146]), .Q(MemoryLatch[146]));
	LATQ_X1M_A12TR MemoryLatch_reg_147(.D(GDIN), .G(DGWCLK[147]), .Q(MemoryLatch[147]));
	LATQ_X1M_A12TR MemoryLatch_reg_148(.D(GDIN), .G(DGWCLK[148]), .Q(MemoryLatch[148]));
	LATQ_X1M_A12TR MemoryLatch_reg_149(.D(GDIN), .G(DGWCLK[149]), .Q(MemoryLatch[149]));
	LATQ_X1M_A12TR MemoryLatch_reg_15(.D(GDIN), .G(DGWCLK[15]), .Q(MemoryLatch[15]));
	LATQ_X1M_A12TR MemoryLatch_reg_150(.D(GDIN), .G(DGWCLK[150]), .Q(MemoryLatch[150]));
	LATQ_X1M_A12TR MemoryLatch_reg_151(.D(GDIN), .G(DGWCLK[151]), .Q(MemoryLatch[151]));
	LATQ_X1M_A12TR MemoryLatch_reg_152(.D(GDIN), .G(DGWCLK[152]), .Q(MemoryLatch[152]));
	LATQ_X1M_A12TR MemoryLatch_reg_153(.D(GDIN), .G(DGWCLK[153]), .Q(MemoryLatch[153]));
	LATQ_X1M_A12TR MemoryLatch_reg_154(.D(GDIN), .G(DGWCLK[154]), .Q(MemoryLatch[154]));
	LATQ_X1M_A12TR MemoryLatch_reg_155(.D(GDIN), .G(DGWCLK[155]), .Q(MemoryLatch[155]));
	LATQ_X1M_A12TR MemoryLatch_reg_156(.D(GDIN), .G(DGWCLK[156]), .Q(MemoryLatch[156]));
	LATQ_X1M_A12TR MemoryLatch_reg_157(.D(GDIN), .G(DGWCLK[157]), .Q(MemoryLatch[157]));
	LATQ_X1M_A12TR MemoryLatch_reg_158(.D(GDIN), .G(DGWCLK[158]), .Q(MemoryLatch[158]));
	LATQ_X1M_A12TR MemoryLatch_reg_159(.D(GDIN), .G(DGWCLK[159]), .Q(MemoryLatch[159]));
	LATQ_X1M_A12TR MemoryLatch_reg_16(.D(GDIN), .G(DGWCLK[16]), .Q(MemoryLatch[16]));
	LATQ_X1M_A12TR MemoryLatch_reg_160(.D(GDIN), .G(DGWCLK[160]), .Q(MemoryLatch[160]));
	LATQ_X1M_A12TR MemoryLatch_reg_161(.D(GDIN), .G(DGWCLK[161]), .Q(MemoryLatch[161]));
	LATQ_X1M_A12TR MemoryLatch_reg_162(.D(GDIN), .G(DGWCLK[162]), .Q(MemoryLatch[162]));
	LATQ_X1M_A12TR MemoryLatch_reg_163(.D(GDIN), .G(DGWCLK[163]), .Q(MemoryLatch[163]));
	LATQ_X1M_A12TR MemoryLatch_reg_164(.D(GDIN), .G(DGWCLK[164]), .Q(MemoryLatch[164]));
	LATQ_X1M_A12TR MemoryLatch_reg_165(.D(GDIN), .G(DGWCLK[165]), .Q(MemoryLatch[165]));
	LATQ_X1M_A12TR MemoryLatch_reg_166(.D(GDIN), .G(DGWCLK[166]), .Q(MemoryLatch[166]));
	LATQ_X1M_A12TR MemoryLatch_reg_167(.D(GDIN), .G(DGWCLK[167]), .Q(MemoryLatch[167]));
	LATQ_X1M_A12TR MemoryLatch_reg_168(.D(GDIN), .G(DGWCLK[168]), .Q(MemoryLatch[168]));
	LATQ_X1M_A12TR MemoryLatch_reg_169(.D(GDIN), .G(DGWCLK[169]), .Q(MemoryLatch[169]));
	LATQ_X1M_A12TR MemoryLatch_reg_17(.D(GDIN), .G(DGWCLK[17]), .Q(MemoryLatch[17]));
	LATQ_X1M_A12TR MemoryLatch_reg_170(.D(GDIN), .G(DGWCLK[170]), .Q(MemoryLatch[170]));
	LATQ_X1M_A12TR MemoryLatch_reg_171(.D(GDIN), .G(DGWCLK[171]), .Q(MemoryLatch[171]));
	LATQ_X1M_A12TR MemoryLatch_reg_172(.D(GDIN), .G(DGWCLK[172]), .Q(MemoryLatch[172]));
	LATQ_X1M_A12TR MemoryLatch_reg_173(.D(GDIN), .G(DGWCLK[173]), .Q(MemoryLatch[173]));
	LATQ_X1M_A12TR MemoryLatch_reg_174(.D(GDIN), .G(DGWCLK[174]), .Q(MemoryLatch[174]));
	LATQ_X1M_A12TR MemoryLatch_reg_175(.D(GDIN), .G(DGWCLK[175]), .Q(MemoryLatch[175]));
	LATQ_X1M_A12TR MemoryLatch_reg_176(.D(GDIN), .G(DGWCLK[176]), .Q(MemoryLatch[176]));
	LATQ_X1M_A12TR MemoryLatch_reg_177(.D(GDIN), .G(DGWCLK[177]), .Q(MemoryLatch[177]));
	LATQ_X1M_A12TR MemoryLatch_reg_178(.D(GDIN), .G(DGWCLK[178]), .Q(MemoryLatch[178]));
	LATQ_X1M_A12TR MemoryLatch_reg_179(.D(GDIN), .G(DGWCLK[179]), .Q(MemoryLatch[179]));
	LATQ_X1M_A12TR MemoryLatch_reg_18(.D(GDIN), .G(DGWCLK[18]), .Q(MemoryLatch[18]));
	LATQ_X1M_A12TR MemoryLatch_reg_180(.D(GDIN), .G(DGWCLK[180]), .Q(MemoryLatch[180]));
	LATQ_X1M_A12TR MemoryLatch_reg_181(.D(GDIN), .G(DGWCLK[181]), .Q(MemoryLatch[181]));
	LATQ_X1M_A12TR MemoryLatch_reg_182(.D(GDIN), .G(DGWCLK[182]), .Q(MemoryLatch[182]));
	LATQ_X1M_A12TR MemoryLatch_reg_183(.D(GDIN), .G(DGWCLK[183]), .Q(MemoryLatch[183]));
	LATQ_X1M_A12TR MemoryLatch_reg_184(.D(GDIN), .G(DGWCLK[184]), .Q(MemoryLatch[184]));
	LATQ_X1M_A12TR MemoryLatch_reg_185(.D(GDIN), .G(DGWCLK[185]), .Q(MemoryLatch[185]));
	LATQ_X1M_A12TR MemoryLatch_reg_186(.D(GDIN), .G(DGWCLK[186]), .Q(MemoryLatch[186]));
	LATQ_X1M_A12TR MemoryLatch_reg_187(.D(GDIN), .G(DGWCLK[187]), .Q(MemoryLatch[187]));
	LATQ_X1M_A12TR MemoryLatch_reg_188(.D(GDIN), .G(DGWCLK[188]), .Q(MemoryLatch[188]));
	LATQ_X1M_A12TR MemoryLatch_reg_189(.D(GDIN), .G(DGWCLK[189]), .Q(MemoryLatch[189]));
	LATQ_X1M_A12TR MemoryLatch_reg_19(.D(GDIN), .G(DGWCLK[19]), .Q(MemoryLatch[19]));
	LATQ_X1M_A12TR MemoryLatch_reg_190(.D(GDIN), .G(DGWCLK[190]), .Q(MemoryLatch[190]));
	LATQ_X1M_A12TR MemoryLatch_reg_191(.D(GDIN), .G(DGWCLK[191]), .Q(MemoryLatch[191]));
	LATQ_X1M_A12TR MemoryLatch_reg_192(.D(GDIN), .G(DGWCLK[192]), .Q(MemoryLatch[192]));
	LATQ_X1M_A12TR MemoryLatch_reg_193(.D(GDIN), .G(DGWCLK[193]), .Q(MemoryLatch[193]));
	LATQ_X1M_A12TR MemoryLatch_reg_194(.D(GDIN), .G(DGWCLK[194]), .Q(MemoryLatch[194]));
	LATQ_X1M_A12TR MemoryLatch_reg_195(.D(GDIN), .G(DGWCLK[195]), .Q(MemoryLatch[195]));
	LATQ_X1M_A12TR MemoryLatch_reg_196(.D(GDIN), .G(DGWCLK[196]), .Q(MemoryLatch[196]));
	LATQ_X1M_A12TR MemoryLatch_reg_197(.D(GDIN), .G(DGWCLK[197]), .Q(MemoryLatch[197]));
	LATQ_X1M_A12TR MemoryLatch_reg_198(.D(GDIN), .G(DGWCLK[198]), .Q(MemoryLatch[198]));
	LATQ_X1M_A12TR MemoryLatch_reg_199(.D(GDIN), .G(DGWCLK[199]), .Q(MemoryLatch[199]));
	LATQ_X1M_A12TR MemoryLatch_reg_2(.D(GDIN), .G(DGWCLK[2]), .Q(MemoryLatch[2]));
	LATQ_X1M_A12TR MemoryLatch_reg_20(.D(GDIN), .G(DGWCLK[20]), .Q(MemoryLatch[20]));
	LATQ_X1M_A12TR MemoryLatch_reg_200(.D(GDIN), .G(DGWCLK[200]), .Q(MemoryLatch[200]));
	LATQ_X1M_A12TR MemoryLatch_reg_201(.D(GDIN), .G(DGWCLK[201]), .Q(MemoryLatch[201]));
	LATQ_X1M_A12TR MemoryLatch_reg_202(.D(GDIN), .G(DGWCLK[202]), .Q(MemoryLatch[202]));
	LATQ_X1M_A12TR MemoryLatch_reg_203(.D(GDIN), .G(DGWCLK[203]), .Q(MemoryLatch[203]));
	LATQ_X1M_A12TR MemoryLatch_reg_204(.D(GDIN), .G(DGWCLK[204]), .Q(MemoryLatch[204]));
	LATQ_X1M_A12TR MemoryLatch_reg_205(.D(GDIN), .G(DGWCLK[205]), .Q(MemoryLatch[205]));
	LATQ_X1M_A12TR MemoryLatch_reg_206(.D(GDIN), .G(DGWCLK[206]), .Q(MemoryLatch[206]));
	LATQ_X1M_A12TR MemoryLatch_reg_207(.D(GDIN), .G(DGWCLK[207]), .Q(MemoryLatch[207]));
	LATQ_X1M_A12TR MemoryLatch_reg_208(.D(GDIN), .G(DGWCLK[208]), .Q(MemoryLatch[208]));
	LATQ_X1M_A12TR MemoryLatch_reg_209(.D(GDIN), .G(DGWCLK[209]), .Q(MemoryLatch[209]));
	LATQ_X1M_A12TR MemoryLatch_reg_21(.D(GDIN), .G(DGWCLK[21]), .Q(MemoryLatch[21]));
	LATQ_X1M_A12TR MemoryLatch_reg_210(.D(GDIN), .G(DGWCLK[210]), .Q(MemoryLatch[210]));
	LATQ_X1M_A12TR MemoryLatch_reg_211(.D(GDIN), .G(DGWCLK[211]), .Q(MemoryLatch[211]));
	LATQ_X1M_A12TR MemoryLatch_reg_212(.D(GDIN), .G(DGWCLK[212]), .Q(MemoryLatch[212]));
	LATQ_X1M_A12TR MemoryLatch_reg_213(.D(GDIN), .G(DGWCLK[213]), .Q(MemoryLatch[213]));
	LATQ_X1M_A12TR MemoryLatch_reg_214(.D(GDIN), .G(DGWCLK[214]), .Q(MemoryLatch[214]));
	LATQ_X1M_A12TR MemoryLatch_reg_215(.D(GDIN), .G(DGWCLK[215]), .Q(MemoryLatch[215]));
	LATQ_X1M_A12TR MemoryLatch_reg_216(.D(GDIN), .G(DGWCLK[216]), .Q(MemoryLatch[216]));
	LATQ_X1M_A12TR MemoryLatch_reg_217(.D(GDIN), .G(DGWCLK[217]), .Q(MemoryLatch[217]));
	LATQ_X1M_A12TR MemoryLatch_reg_218(.D(GDIN), .G(DGWCLK[218]), .Q(MemoryLatch[218]));
	LATQ_X1M_A12TR MemoryLatch_reg_219(.D(GDIN), .G(DGWCLK[219]), .Q(MemoryLatch[219]));
	LATQ_X1M_A12TR MemoryLatch_reg_22(.D(GDIN), .G(DGWCLK[22]), .Q(MemoryLatch[22]));
	LATQ_X1M_A12TR MemoryLatch_reg_220(.D(GDIN), .G(DGWCLK[220]), .Q(MemoryLatch[220]));
	LATQ_X1M_A12TR MemoryLatch_reg_221(.D(GDIN), .G(DGWCLK[221]), .Q(MemoryLatch[221]));
	LATQ_X1M_A12TR MemoryLatch_reg_222(.D(GDIN), .G(DGWCLK[222]), .Q(MemoryLatch[222]));
	LATQ_X1M_A12TR MemoryLatch_reg_223(.D(GDIN), .G(DGWCLK[223]), .Q(MemoryLatch[223]));
	LATQ_X1M_A12TR MemoryLatch_reg_224(.D(GDIN), .G(DGWCLK[224]), .Q(MemoryLatch[224]));
	LATQ_X1M_A12TR MemoryLatch_reg_225(.D(GDIN), .G(DGWCLK[225]), .Q(MemoryLatch[225]));
	LATQ_X1M_A12TR MemoryLatch_reg_226(.D(GDIN), .G(DGWCLK[226]), .Q(MemoryLatch[226]));
	LATQ_X1M_A12TR MemoryLatch_reg_227(.D(GDIN), .G(DGWCLK[227]), .Q(MemoryLatch[227]));
	LATQ_X1M_A12TR MemoryLatch_reg_228(.D(GDIN), .G(DGWCLK[228]), .Q(MemoryLatch[228]));
	LATQ_X1M_A12TR MemoryLatch_reg_229(.D(GDIN), .G(DGWCLK[229]), .Q(MemoryLatch[229]));
	LATQ_X1M_A12TR MemoryLatch_reg_23(.D(GDIN), .G(DGWCLK[23]), .Q(MemoryLatch[23]));
	LATQ_X1M_A12TR MemoryLatch_reg_230(.D(GDIN), .G(DGWCLK[230]), .Q(MemoryLatch[230]));
	LATQ_X1M_A12TR MemoryLatch_reg_231(.D(GDIN), .G(DGWCLK[231]), .Q(MemoryLatch[231]));
	LATQ_X1M_A12TR MemoryLatch_reg_232(.D(GDIN), .G(DGWCLK[232]), .Q(MemoryLatch[232]));
	LATQ_X1M_A12TR MemoryLatch_reg_233(.D(GDIN), .G(DGWCLK[233]), .Q(MemoryLatch[233]));
	LATQ_X1M_A12TR MemoryLatch_reg_234(.D(GDIN), .G(DGWCLK[234]), .Q(MemoryLatch[234]));
	LATQ_X1M_A12TR MemoryLatch_reg_235(.D(GDIN), .G(DGWCLK[235]), .Q(MemoryLatch[235]));
	LATQ_X1M_A12TR MemoryLatch_reg_236(.D(GDIN), .G(DGWCLK[236]), .Q(MemoryLatch[236]));
	LATQ_X1M_A12TR MemoryLatch_reg_237(.D(GDIN), .G(DGWCLK[237]), .Q(MemoryLatch[237]));
	LATQ_X1M_A12TR MemoryLatch_reg_238(.D(GDIN), .G(DGWCLK[238]), .Q(MemoryLatch[238]));
	LATQ_X1M_A12TR MemoryLatch_reg_239(.D(GDIN), .G(DGWCLK[239]), .Q(MemoryLatch[239]));
	LATQ_X1M_A12TR MemoryLatch_reg_24(.D(GDIN), .G(DGWCLK[24]), .Q(MemoryLatch[24]));
	LATQ_X1M_A12TR MemoryLatch_reg_240(.D(GDIN), .G(DGWCLK[240]), .Q(MemoryLatch[240]));
	LATQ_X1M_A12TR MemoryLatch_reg_241(.D(GDIN), .G(DGWCLK[241]), .Q(MemoryLatch[241]));
	LATQ_X1M_A12TR MemoryLatch_reg_242(.D(GDIN), .G(DGWCLK[242]), .Q(MemoryLatch[242]));
	LATQ_X1M_A12TR MemoryLatch_reg_243(.D(GDIN), .G(DGWCLK[243]), .Q(MemoryLatch[243]));
	LATQ_X1M_A12TR MemoryLatch_reg_244(.D(GDIN), .G(DGWCLK[244]), .Q(MemoryLatch[244]));
	LATQ_X1M_A12TR MemoryLatch_reg_245(.D(GDIN), .G(DGWCLK[245]), .Q(MemoryLatch[245]));
	LATQ_X1M_A12TR MemoryLatch_reg_246(.D(GDIN), .G(DGWCLK[246]), .Q(MemoryLatch[246]));
	LATQ_X1M_A12TR MemoryLatch_reg_247(.D(GDIN), .G(DGWCLK[247]), .Q(MemoryLatch[247]));
	LATQ_X1M_A12TR MemoryLatch_reg_248(.D(GDIN), .G(DGWCLK[248]), .Q(MemoryLatch[248]));
	LATQ_X1M_A12TR MemoryLatch_reg_249(.D(GDIN), .G(DGWCLK[249]), .Q(MemoryLatch[249]));
	LATQ_X1M_A12TR MemoryLatch_reg_25(.D(GDIN), .G(DGWCLK[25]), .Q(MemoryLatch[25]));
	LATQ_X1M_A12TR MemoryLatch_reg_250(.D(GDIN), .G(DGWCLK[250]), .Q(MemoryLatch[250]));
	LATQ_X1M_A12TR MemoryLatch_reg_251(.D(GDIN), .G(DGWCLK[251]), .Q(MemoryLatch[251]));
	LATQ_X1M_A12TR MemoryLatch_reg_252(.D(GDIN), .G(DGWCLK[252]), .Q(MemoryLatch[252]));
	LATQ_X1M_A12TR MemoryLatch_reg_253(.D(GDIN), .G(DGWCLK[253]), .Q(MemoryLatch[253]));
	LATQ_X1M_A12TR MemoryLatch_reg_254(.D(GDIN), .G(DGWCLK[254]), .Q(MemoryLatch[254]));
	LATQ_X1M_A12TR MemoryLatch_reg_255(.D(GDIN), .G(DGWCLK[255]), .Q(MemoryLatch[255]));
	LATQ_X1M_A12TR MemoryLatch_reg_26(.D(GDIN), .G(DGWCLK[26]), .Q(MemoryLatch[26]));
	LATQ_X1M_A12TR MemoryLatch_reg_27(.D(GDIN), .G(DGWCLK[27]), .Q(MemoryLatch[27]));
	LATQ_X1M_A12TR MemoryLatch_reg_28(.D(GDIN), .G(DGWCLK[28]), .Q(MemoryLatch[28]));
	LATQ_X1M_A12TR MemoryLatch_reg_29(.D(GDIN), .G(DGWCLK[29]), .Q(MemoryLatch[29]));
	LATQ_X1M_A12TR MemoryLatch_reg_3(.D(GDIN), .G(DGWCLK[3]), .Q(MemoryLatch[3]));
	LATQ_X1M_A12TR MemoryLatch_reg_30(.D(GDIN), .G(DGWCLK[30]), .Q(MemoryLatch[30]));
	LATQ_X1M_A12TR MemoryLatch_reg_31(.D(GDIN), .G(DGWCLK[31]), .Q(MemoryLatch[31]));
	LATQ_X1M_A12TR MemoryLatch_reg_32(.D(GDIN), .G(DGWCLK[32]), .Q(MemoryLatch[32]));
	LATQ_X1M_A12TR MemoryLatch_reg_33(.D(GDIN), .G(DGWCLK[33]), .Q(MemoryLatch[33]));
	LATQ_X1M_A12TR MemoryLatch_reg_34(.D(GDIN), .G(DGWCLK[34]), .Q(MemoryLatch[34]));
	LATQ_X1M_A12TR MemoryLatch_reg_35(.D(GDIN), .G(DGWCLK[35]), .Q(MemoryLatch[35]));
	LATQ_X1M_A12TR MemoryLatch_reg_36(.D(GDIN), .G(DGWCLK[36]), .Q(MemoryLatch[36]));
	LATQ_X1M_A12TR MemoryLatch_reg_37(.D(GDIN), .G(DGWCLK[37]), .Q(MemoryLatch[37]));
	LATQ_X1M_A12TR MemoryLatch_reg_38(.D(GDIN), .G(DGWCLK[38]), .Q(MemoryLatch[38]));
	LATQ_X1M_A12TR MemoryLatch_reg_39(.D(GDIN), .G(DGWCLK[39]), .Q(MemoryLatch[39]));
	LATQ_X1M_A12TR MemoryLatch_reg_4(.D(GDIN), .G(DGWCLK[4]), .Q(MemoryLatch[4]));
	LATQ_X1M_A12TR MemoryLatch_reg_40(.D(GDIN), .G(DGWCLK[40]), .Q(MemoryLatch[40]));
	LATQ_X1M_A12TR MemoryLatch_reg_41(.D(GDIN), .G(DGWCLK[41]), .Q(MemoryLatch[41]));
	LATQ_X1M_A12TR MemoryLatch_reg_42(.D(GDIN), .G(DGWCLK[42]), .Q(MemoryLatch[42]));
	LATQ_X1M_A12TR MemoryLatch_reg_43(.D(GDIN), .G(DGWCLK[43]), .Q(MemoryLatch[43]));
	LATQ_X1M_A12TR MemoryLatch_reg_44(.D(GDIN), .G(DGWCLK[44]), .Q(MemoryLatch[44]));
	LATQ_X1M_A12TR MemoryLatch_reg_45(.D(GDIN), .G(DGWCLK[45]), .Q(MemoryLatch[45]));
	LATQ_X1M_A12TR MemoryLatch_reg_46(.D(GDIN), .G(DGWCLK[46]), .Q(MemoryLatch[46]));
	LATQ_X1M_A12TR MemoryLatch_reg_47(.D(GDIN), .G(DGWCLK[47]), .Q(MemoryLatch[47]));
	LATQ_X1M_A12TR MemoryLatch_reg_48(.D(GDIN), .G(DGWCLK[48]), .Q(MemoryLatch[48]));
	LATQ_X1M_A12TR MemoryLatch_reg_49(.D(GDIN), .G(DGWCLK[49]), .Q(MemoryLatch[49]));
	LATQ_X1M_A12TR MemoryLatch_reg_5(.D(GDIN), .G(DGWCLK[5]), .Q(MemoryLatch[5]));
	LATQ_X1M_A12TR MemoryLatch_reg_50(.D(GDIN), .G(DGWCLK[50]), .Q(MemoryLatch[50]));
	LATQ_X1M_A12TR MemoryLatch_reg_51(.D(GDIN), .G(DGWCLK[51]), .Q(MemoryLatch[51]));
	LATQ_X1M_A12TR MemoryLatch_reg_52(.D(GDIN), .G(DGWCLK[52]), .Q(MemoryLatch[52]));
	LATQ_X1M_A12TR MemoryLatch_reg_53(.D(GDIN), .G(DGWCLK[53]), .Q(MemoryLatch[53]));
	LATQ_X1M_A12TR MemoryLatch_reg_54(.D(GDIN), .G(DGWCLK[54]), .Q(MemoryLatch[54]));
	LATQ_X1M_A12TR MemoryLatch_reg_55(.D(GDIN), .G(DGWCLK[55]), .Q(MemoryLatch[55]));
	LATQ_X1M_A12TR MemoryLatch_reg_56(.D(GDIN), .G(DGWCLK[56]), .Q(MemoryLatch[56]));
	LATQ_X1M_A12TR MemoryLatch_reg_57(.D(GDIN), .G(DGWCLK[57]), .Q(MemoryLatch[57]));
	LATQ_X1M_A12TR MemoryLatch_reg_58(.D(GDIN), .G(DGWCLK[58]), .Q(MemoryLatch[58]));
	LATQ_X1M_A12TR MemoryLatch_reg_59(.D(GDIN), .G(DGWCLK[59]), .Q(MemoryLatch[59]));
	LATQ_X1M_A12TR MemoryLatch_reg_6(.D(GDIN), .G(DGWCLK[6]), .Q(MemoryLatch[6]));
	LATQ_X1M_A12TR MemoryLatch_reg_60(.D(GDIN), .G(DGWCLK[60]), .Q(MemoryLatch[60]));
	LATQ_X1M_A12TR MemoryLatch_reg_61(.D(GDIN), .G(DGWCLK[61]), .Q(MemoryLatch[61]));
	LATQ_X1M_A12TR MemoryLatch_reg_62(.D(GDIN), .G(DGWCLK[62]), .Q(MemoryLatch[62]));
	LATQ_X1M_A12TR MemoryLatch_reg_63(.D(GDIN), .G(DGWCLK[63]), .Q(MemoryLatch[63]));
	LATQ_X1M_A12TR MemoryLatch_reg_64(.D(GDIN), .G(DGWCLK[64]), .Q(MemoryLatch[64]));
	LATQ_X1M_A12TR MemoryLatch_reg_65(.D(GDIN), .G(DGWCLK[65]), .Q(MemoryLatch[65]));
	LATQ_X1M_A12TR MemoryLatch_reg_66(.D(GDIN), .G(DGWCLK[66]), .Q(MemoryLatch[66]));
	LATQ_X1M_A12TR MemoryLatch_reg_67(.D(GDIN), .G(DGWCLK[67]), .Q(MemoryLatch[67]));
	LATQ_X1M_A12TR MemoryLatch_reg_68(.D(GDIN), .G(DGWCLK[68]), .Q(MemoryLatch[68]));
	LATQ_X1M_A12TR MemoryLatch_reg_69(.D(GDIN), .G(DGWCLK[69]), .Q(MemoryLatch[69]));
	LATQ_X1M_A12TR MemoryLatch_reg_7(.D(GDIN), .G(DGWCLK[7]), .Q(MemoryLatch[7]));
	LATQ_X1M_A12TR MemoryLatch_reg_70(.D(GDIN), .G(DGWCLK[70]), .Q(MemoryLatch[70]));
	LATQ_X1M_A12TR MemoryLatch_reg_71(.D(GDIN), .G(DGWCLK[71]), .Q(MemoryLatch[71]));
	LATQ_X1M_A12TR MemoryLatch_reg_72(.D(GDIN), .G(DGWCLK[72]), .Q(MemoryLatch[72]));
	LATQ_X1M_A12TR MemoryLatch_reg_73(.D(GDIN), .G(DGWCLK[73]), .Q(MemoryLatch[73]));
	LATQ_X1M_A12TR MemoryLatch_reg_74(.D(GDIN), .G(DGWCLK[74]), .Q(MemoryLatch[74]));
	LATQ_X1M_A12TR MemoryLatch_reg_75(.D(GDIN), .G(DGWCLK[75]), .Q(MemoryLatch[75]));
	LATQ_X1M_A12TR MemoryLatch_reg_76(.D(GDIN), .G(DGWCLK[76]), .Q(MemoryLatch[76]));
	LATQ_X1M_A12TR MemoryLatch_reg_77(.D(GDIN), .G(DGWCLK[77]), .Q(MemoryLatch[77]));
	LATQ_X1M_A12TR MemoryLatch_reg_78(.D(GDIN), .G(DGWCLK[78]), .Q(MemoryLatch[78]));
	LATQ_X1M_A12TR MemoryLatch_reg_79(.D(GDIN), .G(DGWCLK[79]), .Q(MemoryLatch[79]));
	LATQ_X1M_A12TR MemoryLatch_reg_8(.D(GDIN), .G(DGWCLK[8]), .Q(MemoryLatch[8]));
	LATQ_X1M_A12TR MemoryLatch_reg_80(.D(GDIN), .G(DGWCLK[80]), .Q(MemoryLatch[80]));
	LATQ_X1M_A12TR MemoryLatch_reg_81(.D(GDIN), .G(DGWCLK[81]), .Q(MemoryLatch[81]));
	LATQ_X1M_A12TR MemoryLatch_reg_82(.D(GDIN), .G(DGWCLK[82]), .Q(MemoryLatch[82]));
	LATQ_X1M_A12TR MemoryLatch_reg_83(.D(GDIN), .G(DGWCLK[83]), .Q(MemoryLatch[83]));
	LATQ_X1M_A12TR MemoryLatch_reg_84(.D(GDIN), .G(DGWCLK[84]), .Q(MemoryLatch[84]));
	LATQ_X1M_A12TR MemoryLatch_reg_85(.D(GDIN), .G(DGWCLK[85]), .Q(MemoryLatch[85]));
	LATQ_X1M_A12TR MemoryLatch_reg_86(.D(GDIN), .G(DGWCLK[86]), .Q(MemoryLatch[86]));
	LATQ_X1M_A12TR MemoryLatch_reg_87(.D(GDIN), .G(DGWCLK[87]), .Q(MemoryLatch[87]));
	LATQ_X1M_A12TR MemoryLatch_reg_88(.D(GDIN), .G(DGWCLK[88]), .Q(MemoryLatch[88]));
	LATQ_X1M_A12TR MemoryLatch_reg_89(.D(GDIN), .G(DGWCLK[89]), .Q(MemoryLatch[89]));
	LATQ_X1M_A12TR MemoryLatch_reg_9(.D(GDIN), .G(DGWCLK[9]), .Q(MemoryLatch[9]));
	LATQ_X1M_A12TR MemoryLatch_reg_90(.D(GDIN), .G(DGWCLK[90]), .Q(MemoryLatch[90]));
	LATQ_X1M_A12TR MemoryLatch_reg_91(.D(GDIN), .G(DGWCLK[91]), .Q(MemoryLatch[91]));
	LATQ_X1M_A12TR MemoryLatch_reg_92(.D(GDIN), .G(DGWCLK[92]), .Q(MemoryLatch[92]));
	LATQ_X1M_A12TR MemoryLatch_reg_93(.D(GDIN), .G(DGWCLK[93]), .Q(MemoryLatch[93]));
	LATQ_X1M_A12TR MemoryLatch_reg_94(.D(GDIN), .G(DGWCLK[94]), .Q(MemoryLatch[94]));
	LATQ_X1M_A12TR MemoryLatch_reg_95(.D(GDIN), .G(DGWCLK[95]), .Q(MemoryLatch[95]));
	LATQ_X1M_A12TR MemoryLatch_reg_96(.D(GDIN), .G(DGWCLK[96]), .Q(MemoryLatch[96]));
	LATQ_X1M_A12TR MemoryLatch_reg_97(.D(GDIN), .G(DGWCLK[97]), .Q(MemoryLatch[97]));
	LATQ_X1M_A12TR MemoryLatch_reg_98(.D(GDIN), .G(DGWCLK[98]), .Q(MemoryLatch[98]));
	LATQ_X1M_A12TR MemoryLatch_reg_99(.D(GDIN), .G(DGWCLK[99]), .Q(MemoryLatch[99]));
	read_mux read_mux(.DOUT(DOUT), .MemoryLatch({MemoryLatch[255:0]}), .RWL({RWL[255:0]}));

endmodule
